-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity mul_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end mul_0CLK_64d180f1;
architecture arch of mul_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1969_c6_4f75]
signal BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1969_c2_7d0a]
signal n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1969_c2_7d0a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1969_c2_7d0a]
signal result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1969_c2_7d0a]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1969_c2_7d0a]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1969_c2_7d0a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1969_c2_7d0a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1969_c2_7d0a]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1969_c2_7d0a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1969_c2_7d0a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1969_c2_7d0a]
signal t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1982_c11_c983]
signal BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1982_c7_dac1]
signal n8_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1982_c7_dac1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1982_c7_dac1]
signal result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1982_c7_dac1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1982_c7_dac1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1982_c7_dac1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1982_c7_dac1]
signal t8_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1985_c11_6c53]
signal BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1985_c7_599f]
signal n8_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1985_c7_599f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1985_c7_599f]
signal result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1985_c7_599f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1985_c7_599f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1985_c7_599f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1985_c7_599f]
signal t8_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1988_c11_e782]
signal BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1988_c7_5236]
signal n8_MUX_uxn_opcodes_h_l1988_c7_5236_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1988_c7_5236_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1988_c7_5236]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1988_c7_5236]
signal result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1988_c7_5236]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1988_c7_5236]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1988_c7_5236]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1990_c30_8cd0]
signal sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_return_output : signed(3 downto 0);

-- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1993_c21_d83c]
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_left : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_right : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_return_output : unsigned(15 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_b856( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75
BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_left,
BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_right,
BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output);

-- n8_MUX_uxn_opcodes_h_l1969_c2_7d0a
n8_MUX_uxn_opcodes_h_l1969_c2_7d0a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond,
n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue,
n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse,
n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a
result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a
result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a
result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a
result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a
result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a
result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output);

-- t8_MUX_uxn_opcodes_h_l1969_c2_7d0a
t8_MUX_uxn_opcodes_h_l1969_c2_7d0a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond,
t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue,
t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse,
t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983
BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_left,
BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_right,
BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_return_output);

-- n8_MUX_uxn_opcodes_h_l1982_c7_dac1
n8_MUX_uxn_opcodes_h_l1982_c7_dac1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1982_c7_dac1_cond,
n8_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue,
n8_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse,
n8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1
result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_cond,
result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1
result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1
result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1
result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output);

-- t8_MUX_uxn_opcodes_h_l1982_c7_dac1
t8_MUX_uxn_opcodes_h_l1982_c7_dac1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1982_c7_dac1_cond,
t8_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue,
t8_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse,
t8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53
BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_left,
BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_right,
BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_return_output);

-- n8_MUX_uxn_opcodes_h_l1985_c7_599f
n8_MUX_uxn_opcodes_h_l1985_c7_599f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1985_c7_599f_cond,
n8_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue,
n8_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse,
n8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f
result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f
result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f
result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_return_output);

-- t8_MUX_uxn_opcodes_h_l1985_c7_599f
t8_MUX_uxn_opcodes_h_l1985_c7_599f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1985_c7_599f_cond,
t8_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue,
t8_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse,
t8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782
BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_left,
BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_right,
BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_return_output);

-- n8_MUX_uxn_opcodes_h_l1988_c7_5236
n8_MUX_uxn_opcodes_h_l1988_c7_5236 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1988_c7_5236_cond,
n8_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue,
n8_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse,
n8_MUX_uxn_opcodes_h_l1988_c7_5236_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236
result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_cond,
result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236
result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236
result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236
result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0
sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_ins,
sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_x,
sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_y,
sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_return_output);

-- BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c : entity work.BIN_OP_INFERRED_MULT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_left,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_right,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output,
 n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
 t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_return_output,
 n8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output,
 t8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_return_output,
 n8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_return_output,
 t8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_return_output,
 n8_MUX_uxn_opcodes_h_l1988_c7_5236_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_return_output,
 sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_return_output,
 BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1979_c3_5d82 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1974_c3_830a : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1983_c3_817b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1982_c7_dac1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1988_c7_5236_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1985_c7_599f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1988_c7_5236_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1992_c3_7d61 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l1993_c3_b2fa : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1985_l1969_l1988_l1982_DUPLICATE_5ce1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_0b35_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_a421_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_bd85_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1985_l1988_DUPLICATE_d0d0_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1997_l1965_DUPLICATE_a49e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1974_c3_830a := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1974_c3_830a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_right := to_unsigned(2, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1992_c3_7d61 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1992_c3_7d61;
     VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1983_c3_817b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1983_c3_817b;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1979_c3_5d82 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1979_c3_5d82;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_left := VAR_phase;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1969_c6_4f75] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_left;
     BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output := BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output;

     -- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1993_c21_d83c] LATENCY=0
     -- Inputs
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_left <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_left;
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_right <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_right;
     -- Outputs
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_return_output := BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1985_l1969_l1988_l1982_DUPLICATE_5ce1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1985_l1969_l1988_l1982_DUPLICATE_5ce1_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1982_c11_c983] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_left;
     BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_return_output := BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1985_c11_6c53] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_left;
     BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_return_output := BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_bd85 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_bd85_return_output := result.is_opc_done;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1969_c2_7d0a_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_0b35 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_0b35_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1985_l1988_DUPLICATE_d0d0 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1985_l1988_DUPLICATE_d0d0_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1988_c11_e782] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_left;
     BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_return_output := BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1990_c30_8cd0] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_ins;
     sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_x;
     sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_return_output := sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1969_c2_7d0a_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_a421 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_a421_return_output := result.sp_relative_shift;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1969_c2_7d0a_return_output := result.is_vram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1969_c2_7d0a_return_output := result.is_pc_updated;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_4f75_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1982_c7_dac1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1982_c7_dac1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_c983_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1985_c7_599f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1985_c7_599f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_6c53_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1988_c7_5236_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_e782_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l1993_c3_b2fa := resize(VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_d83c_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_a421_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_a421_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_a421_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_bd85_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_bd85_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_bd85_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_0b35_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_0b35_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1985_l1988_l1982_DUPLICATE_0b35_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1985_l1988_DUPLICATE_d0d0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1985_l1988_DUPLICATE_d0d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1985_l1969_l1988_l1982_DUPLICATE_5ce1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1985_l1969_l1988_l1982_DUPLICATE_5ce1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1985_l1969_l1988_l1982_DUPLICATE_5ce1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1985_l1969_l1988_l1982_DUPLICATE_5ce1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1969_c2_7d0a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1969_c2_7d0a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1969_c2_7d0a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1969_c2_7d0a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_8cd0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue := VAR_result_u8_value_uxn_opcodes_h_l1993_c3_b2fa;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1988_c7_5236] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_return_output;

     -- n8_MUX[uxn_opcodes_h_l1988_c7_5236] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1988_c7_5236_cond <= VAR_n8_MUX_uxn_opcodes_h_l1988_c7_5236_cond;
     n8_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue;
     n8_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1988_c7_5236_return_output := n8_MUX_uxn_opcodes_h_l1988_c7_5236_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1988_c7_5236] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1988_c7_5236] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1988_c7_5236] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_return_output := result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1988_c7_5236] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_return_output;

     -- t8_MUX[uxn_opcodes_h_l1985_c7_599f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1985_c7_599f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1985_c7_599f_cond;
     t8_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue;
     t8_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output := t8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1988_c7_5236_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_5236_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_5236_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_5236_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_5236_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_5236_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1985_c7_599f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1985_c7_599f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;

     -- n8_MUX[uxn_opcodes_h_l1985_c7_599f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1985_c7_599f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1985_c7_599f_cond;
     n8_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue;
     n8_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output := n8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1982_c7_dac1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1982_c7_dac1_cond <= VAR_t8_MUX_uxn_opcodes_h_l1982_c7_dac1_cond;
     t8_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue;
     t8_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output := t8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1985_c7_599f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1985_c7_599f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1985_c7_599f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_599f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1982_c7_dac1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output := result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1982_c7_dac1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;

     -- t8_MUX[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond;
     t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue;
     t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output := t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1982_c7_dac1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1982_c7_dac1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;

     -- n8_MUX[uxn_opcodes_h_l1982_c7_dac1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1982_c7_dac1_cond <= VAR_n8_MUX_uxn_opcodes_h_l1982_c7_dac1_cond;
     n8_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue;
     n8_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output := n8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1982_c7_dac1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_dac1_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output;

     -- n8_MUX[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond <= VAR_n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond;
     n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue;
     n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output := n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1969_c2_7d0a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1997_l1965_DUPLICATE_a49e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1997_l1965_DUPLICATE_a49e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_b856(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_7d0a_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1997_l1965_DUPLICATE_a49e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1997_l1965_DUPLICATE_a49e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
