-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity eor_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor_0CLK_bacf6a1d;
architecture arch of eor_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1035_c6_f47d]
signal BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1035_c1_51e2]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1035_c2_3520]
signal t8_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1035_c2_3520]
signal n8_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1035_c2_3520]
signal result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1035_c2_3520]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1035_c2_3520]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1035_c2_3520]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1035_c2_3520]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1035_c2_3520]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l1036_c3_debf[uxn_opcodes_h_l1036_c3_debf]
signal printf_uxn_opcodes_h_l1036_c3_debf_uxn_opcodes_h_l1036_c3_debf_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1040_c11_3415]
signal BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1040_c7_1b6b]
signal t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1040_c7_1b6b]
signal n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1040_c7_1b6b]
signal result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1040_c7_1b6b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1040_c7_1b6b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1040_c7_1b6b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1040_c7_1b6b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1040_c7_1b6b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1043_c11_ba93]
signal BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1043_c7_e121]
signal t8_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1043_c7_e121]
signal n8_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1043_c7_e121]
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1043_c7_e121]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1043_c7_e121]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1043_c7_e121]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1043_c7_e121]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1043_c7_e121]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1046_c11_f705]
signal BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1046_c7_c7c2]
signal n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1046_c7_c7c2]
signal result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1046_c7_c7c2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1046_c7_c7c2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1046_c7_c7c2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1046_c7_c7c2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1046_c7_c7c2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1049_c30_c6c0]
signal sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_return_output : signed(3 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1052_c21_4eb8]
signal BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_left : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_right : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1054_c11_61db]
signal BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1054_c7_2dfa]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1054_c7_2dfa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1054_c7_2dfa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d
BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_left,
BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_right,
BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_return_output);

-- t8_MUX_uxn_opcodes_h_l1035_c2_3520
t8_MUX_uxn_opcodes_h_l1035_c2_3520 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1035_c2_3520_cond,
t8_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue,
t8_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse,
t8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output);

-- n8_MUX_uxn_opcodes_h_l1035_c2_3520
n8_MUX_uxn_opcodes_h_l1035_c2_3520 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1035_c2_3520_cond,
n8_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue,
n8_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse,
n8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_cond,
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output);

-- printf_uxn_opcodes_h_l1036_c3_debf_uxn_opcodes_h_l1036_c3_debf
printf_uxn_opcodes_h_l1036_c3_debf_uxn_opcodes_h_l1036_c3_debf : entity work.printf_uxn_opcodes_h_l1036_c3_debf_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1036_c3_debf_uxn_opcodes_h_l1036_c3_debf_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415
BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_left,
BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_right,
BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output);

-- t8_MUX_uxn_opcodes_h_l1040_c7_1b6b
t8_MUX_uxn_opcodes_h_l1040_c7_1b6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond,
t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue,
t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse,
t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output);

-- n8_MUX_uxn_opcodes_h_l1040_c7_1b6b
n8_MUX_uxn_opcodes_h_l1040_c7_1b6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond,
n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue,
n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse,
n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93
BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_left,
BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_right,
BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output);

-- t8_MUX_uxn_opcodes_h_l1043_c7_e121
t8_MUX_uxn_opcodes_h_l1043_c7_e121 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1043_c7_e121_cond,
t8_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue,
t8_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse,
t8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output);

-- n8_MUX_uxn_opcodes_h_l1043_c7_e121
n8_MUX_uxn_opcodes_h_l1043_c7_e121 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1043_c7_e121_cond,
n8_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue,
n8_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse,
n8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_cond,
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705
BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_left,
BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_right,
BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_return_output);

-- n8_MUX_uxn_opcodes_h_l1046_c7_c7c2
n8_MUX_uxn_opcodes_h_l1046_c7_c7c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond,
n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue,
n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse,
n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0
sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_ins,
sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_x,
sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_y,
sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8
BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8 : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_left,
BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_right,
BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db
BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_left,
BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_right,
BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_return_output,
 t8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output,
 n8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output,
 t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output,
 n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output,
 t8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output,
 n8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_return_output,
 n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output,
 sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1037_c3_ba49 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1036_c3_debf_uxn_opcodes_h_l1036_c3_debf_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1041_c3_6c37 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1051_c3_0ce4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_17e0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_ae04_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_b8f4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_a6b9_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1043_l1046_l1040_l1054_DUPLICATE_2c51_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_5286_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1060_l1031_DUPLICATE_b510_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1051_c3_0ce4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1051_c3_0ce4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1037_c3_ba49 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1037_c3_ba49;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1041_c3_6c37 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1041_c3_6c37;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1054_c11_61db] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_left;
     BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_return_output := BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_return_output;

     -- BIN_OP_XOR[uxn_opcodes_h_l1052_c21_4eb8] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_left;
     BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_return_output := BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1046_c11_f705] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_left;
     BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_return_output := BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_ae04 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_ae04_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_17e0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_17e0_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_a6b9 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_a6b9_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l1049_c30_c6c0] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_ins;
     sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_x;
     sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_return_output := sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_b8f4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_b8f4_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1040_c11_3415] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_left;
     BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output := BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1035_c6_f47d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_5286 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_5286_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1043_l1046_l1040_l1054_DUPLICATE_2c51 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1043_l1046_l1040_l1054_DUPLICATE_2c51_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1043_c11_ba93] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_left;
     BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output := BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1035_c2_3520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1035_c2_3520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f47d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_3415_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1043_c7_e121_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1043_c7_e121_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_ba93_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_f705_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_61db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_4eb8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_a6b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_a6b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_a6b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_a6b9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1043_l1046_l1040_l1054_DUPLICATE_2c51_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1043_l1046_l1040_l1054_DUPLICATE_2c51_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1043_l1046_l1040_l1054_DUPLICATE_2c51_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1043_l1046_l1040_l1054_DUPLICATE_2c51_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_ae04_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_ae04_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_ae04_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_ae04_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_b8f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_b8f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_b8f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1043_l1035_l1040_l1054_DUPLICATE_b8f4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_5286_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_5286_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_17e0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_17e0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_17e0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_17e0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_c6c0_return_output;
     -- n8_MUX[uxn_opcodes_h_l1046_c7_c7c2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond <= VAR_n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond;
     n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue;
     n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output := n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1046_c7_c7c2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1035_c1_51e2] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1054_c7_2dfa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1054_c7_2dfa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1046_c7_c7c2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1046_c7_c7c2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;

     -- t8_MUX[uxn_opcodes_h_l1043_c7_e121] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1043_c7_e121_cond <= VAR_t8_MUX_uxn_opcodes_h_l1043_c7_e121_cond;
     t8_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue;
     t8_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output := t8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1054_c7_2dfa] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l1036_c3_debf_uxn_opcodes_h_l1036_c3_debf_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_51e2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_2dfa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1043_c7_e121] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;

     -- t8_MUX[uxn_opcodes_h_l1040_c7_1b6b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond;
     t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue;
     t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output := t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;

     -- printf_uxn_opcodes_h_l1036_c3_debf[uxn_opcodes_h_l1036_c3_debf] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1036_c3_debf_uxn_opcodes_h_l1036_c3_debf_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1036_c3_debf_uxn_opcodes_h_l1036_c3_debf_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1046_c7_c7c2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1046_c7_c7c2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;

     -- n8_MUX[uxn_opcodes_h_l1043_c7_e121] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1043_c7_e121_cond <= VAR_n8_MUX_uxn_opcodes_h_l1043_c7_e121_cond;
     n8_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue;
     n8_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output := n8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1046_c7_c7c2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1043_c7_e121] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1043_c7_e121] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_return_output := result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_c7c2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1040_c7_1b6b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1040_c7_1b6b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1043_c7_e121] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1040_c7_1b6b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1043_c7_e121] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1043_c7_e121] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;

     -- t8_MUX[uxn_opcodes_h_l1035_c2_3520] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1035_c2_3520_cond <= VAR_t8_MUX_uxn_opcodes_h_l1035_c2_3520_cond;
     t8_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue;
     t8_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output := t8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output;

     -- n8_MUX[uxn_opcodes_h_l1040_c7_1b6b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond;
     n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue;
     n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output := n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_e121_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1035_c2_3520] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1035_c2_3520] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_return_output := result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_return_output;

     -- n8_MUX[uxn_opcodes_h_l1035_c2_3520] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1035_c2_3520_cond <= VAR_n8_MUX_uxn_opcodes_h_l1035_c2_3520_cond;
     n8_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue;
     n8_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output := n8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1040_c7_1b6b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1040_c7_1b6b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1040_c7_1b6b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1035_c2_3520] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1035_c2_3520_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_1b6b_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1035_c2_3520] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1035_c2_3520] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1035_c2_3520] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1060_l1031_DUPLICATE_b510 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1060_l1031_DUPLICATE_b510_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_3520_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_3520_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_3520_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_3520_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_3520_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1060_l1031_DUPLICATE_b510_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1060_l1031_DUPLICATE_b510_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
