-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity equ_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_226c8821;
architecture arch of equ_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1162_c6_79b2]
signal BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1162_c2_4851]
signal n8_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1162_c2_4851]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1162_c2_4851]
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1162_c2_4851]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1162_c2_4851]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1162_c2_4851]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1162_c2_4851]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1162_c2_4851]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1162_c2_4851]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1162_c2_4851]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1162_c2_4851]
signal t8_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1175_c11_0867]
signal BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1175_c7_b43e]
signal n8_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1175_c7_b43e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1175_c7_b43e]
signal result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1175_c7_b43e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1175_c7_b43e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1175_c7_b43e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1175_c7_b43e]
signal t8_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1178_c11_b2c4]
signal BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1178_c7_5aed]
signal n8_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1178_c7_5aed]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1178_c7_5aed]
signal result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1178_c7_5aed]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1178_c7_5aed]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1178_c7_5aed]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1178_c7_5aed]
signal t8_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1181_c11_56f6]
signal BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1181_c7_bbbe]
signal n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1181_c7_bbbe]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1181_c7_bbbe]
signal result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1181_c7_bbbe]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1181_c7_bbbe]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1181_c7_bbbe]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1183_c30_3bda]
signal sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1186_c21_c5f4]
signal BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1186_c21_f28d]
signal MUX_uxn_opcodes_h_l1186_c21_f28d_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1186_c21_f28d_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1186_c21_f28d_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1186_c21_f28d_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_b856( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_left,
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_right,
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output);

-- n8_MUX_uxn_opcodes_h_l1162_c2_4851
n8_MUX_uxn_opcodes_h_l1162_c2_4851 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1162_c2_4851_cond,
n8_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue,
n8_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse,
n8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_cond,
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_return_output);

-- t8_MUX_uxn_opcodes_h_l1162_c2_4851
t8_MUX_uxn_opcodes_h_l1162_c2_4851 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1162_c2_4851_cond,
t8_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue,
t8_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse,
t8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867
BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_left,
BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_right,
BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_return_output);

-- n8_MUX_uxn_opcodes_h_l1175_c7_b43e
n8_MUX_uxn_opcodes_h_l1175_c7_b43e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1175_c7_b43e_cond,
n8_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue,
n8_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse,
n8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output);

-- t8_MUX_uxn_opcodes_h_l1175_c7_b43e
t8_MUX_uxn_opcodes_h_l1175_c7_b43e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1175_c7_b43e_cond,
t8_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue,
t8_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse,
t8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4
BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_left,
BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_right,
BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_return_output);

-- n8_MUX_uxn_opcodes_h_l1178_c7_5aed
n8_MUX_uxn_opcodes_h_l1178_c7_5aed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1178_c7_5aed_cond,
n8_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue,
n8_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse,
n8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_cond,
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output);

-- t8_MUX_uxn_opcodes_h_l1178_c7_5aed
t8_MUX_uxn_opcodes_h_l1178_c7_5aed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1178_c7_5aed_cond,
t8_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue,
t8_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse,
t8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6
BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_left,
BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_right,
BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_return_output);

-- n8_MUX_uxn_opcodes_h_l1181_c7_bbbe
n8_MUX_uxn_opcodes_h_l1181_c7_bbbe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond,
n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue,
n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse,
n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond,
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda
sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_ins,
sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_x,
sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_y,
sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4
BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_left,
BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_right,
BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_return_output);

-- MUX_uxn_opcodes_h_l1186_c21_f28d
MUX_uxn_opcodes_h_l1186_c21_f28d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1186_c21_f28d_cond,
MUX_uxn_opcodes_h_l1186_c21_f28d_iftrue,
MUX_uxn_opcodes_h_l1186_c21_f28d_iffalse,
MUX_uxn_opcodes_h_l1186_c21_f28d_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output,
 n8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
 t8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_return_output,
 n8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output,
 t8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_return_output,
 n8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output,
 t8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_return_output,
 n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output,
 sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_return_output,
 MUX_uxn_opcodes_h_l1186_c21_f28d_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1172_c3_ea88 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1167_c3_3484 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1162_c2_4851_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1176_c3_a74c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1175_c7_b43e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5aed_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1185_c3_7840 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1186_c21_f28d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1186_c21_f28d_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1186_c21_f28d_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1186_c21_f28d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1162_l1181_l1178_DUPLICATE_022c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_1a07_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_c599_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_b52e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1181_l1178_DUPLICATE_c7d6_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1190_l1158_DUPLICATE_9705_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1185_c3_7840 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1185_c3_7840;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1176_c3_a74c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1176_c3_a74c;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_right := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_y := resize(to_signed(-1, 2), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1167_c3_3484 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1167_c3_3484;
     VAR_MUX_uxn_opcodes_h_l1186_c21_f28d_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1186_c21_f28d_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1172_c3_ea88 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1172_c3_ea88;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1162_c6_79b2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1186_c21_c5f4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_b52e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_b52e_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1175_c11_0867] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_left;
     BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_return_output := BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1162_l1181_l1178_DUPLICATE_022c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1162_l1181_l1178_DUPLICATE_022c_return_output := result.u8_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1162_c2_4851_return_output := result.is_ram_write;

     -- sp_relative_shift[uxn_opcodes_h_l1183_c30_3bda] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_ins;
     sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_x;
     sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_return_output := sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1162_c2_4851_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1181_c11_56f6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_left;
     BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_return_output := BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_c599 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_c599_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_1a07 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_1a07_return_output := result.is_stack_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1162_c2_4851_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1178_c11_b2c4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1162_c2_4851_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1181_l1178_DUPLICATE_c7d6 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1181_l1178_DUPLICATE_c7d6_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1162_c2_4851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1162_c2_4851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_79b2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1175_c7_b43e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1175_c7_b43e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_0867_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_b2c4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_56f6_return_output;
     VAR_MUX_uxn_opcodes_h_l1186_c21_f28d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_c5f4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_c599_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_c599_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_c599_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_b52e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_b52e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_b52e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_1a07_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_1a07_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1175_l1181_l1178_DUPLICATE_1a07_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1181_l1178_DUPLICATE_c7d6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1181_l1178_DUPLICATE_c7d6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1162_l1181_l1178_DUPLICATE_022c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1162_l1181_l1178_DUPLICATE_022c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1162_l1181_l1178_DUPLICATE_022c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1175_l1162_l1181_l1178_DUPLICATE_022c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1162_c2_4851_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1162_c2_4851_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1162_c2_4851_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1162_c2_4851_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_3bda_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1181_c7_bbbe] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1181_c7_bbbe] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output;

     -- n8_MUX[uxn_opcodes_h_l1181_c7_bbbe] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond <= VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond;
     n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue;
     n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output := n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1181_c7_bbbe] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1181_c7_bbbe] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output;

     -- MUX[uxn_opcodes_h_l1186_c21_f28d] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1186_c21_f28d_cond <= VAR_MUX_uxn_opcodes_h_l1186_c21_f28d_cond;
     MUX_uxn_opcodes_h_l1186_c21_f28d_iftrue <= VAR_MUX_uxn_opcodes_h_l1186_c21_f28d_iftrue;
     MUX_uxn_opcodes_h_l1186_c21_f28d_iffalse <= VAR_MUX_uxn_opcodes_h_l1186_c21_f28d_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1186_c21_f28d_return_output := MUX_uxn_opcodes_h_l1186_c21_f28d_return_output;

     -- t8_MUX[uxn_opcodes_h_l1178_c7_5aed] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1178_c7_5aed_cond <= VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5aed_cond;
     t8_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue;
     t8_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output := t8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue := VAR_MUX_uxn_opcodes_h_l1186_c21_f28d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1178_c7_5aed] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1178_c7_5aed] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1178_c7_5aed] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1178_c7_5aed] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;

     -- t8_MUX[uxn_opcodes_h_l1175_c7_b43e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1175_c7_b43e_cond <= VAR_t8_MUX_uxn_opcodes_h_l1175_c7_b43e_cond;
     t8_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue;
     t8_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output := t8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1181_c7_bbbe] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output := result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output;

     -- n8_MUX[uxn_opcodes_h_l1178_c7_5aed] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1178_c7_5aed_cond <= VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5aed_cond;
     n8_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue;
     n8_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output := n8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_bbbe_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1175_c7_b43e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;

     -- n8_MUX[uxn_opcodes_h_l1175_c7_b43e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1175_c7_b43e_cond <= VAR_n8_MUX_uxn_opcodes_h_l1175_c7_b43e_cond;
     n8_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue;
     n8_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output := n8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1175_c7_b43e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;

     -- t8_MUX[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1162_c2_4851_cond <= VAR_t8_MUX_uxn_opcodes_h_l1162_c2_4851_cond;
     t8_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue;
     t8_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output := t8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1178_c7_5aed] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output := result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1175_c7_b43e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1175_c7_b43e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5aed_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1175_c7_b43e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output;

     -- n8_MUX[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1162_c2_4851_cond <= VAR_n8_MUX_uxn_opcodes_h_l1162_c2_4851_cond;
     n8_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue;
     n8_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output := n8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1162_c2_4851_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_b43e_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1162_c2_4851] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_return_output := result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1190_l1158_DUPLICATE_9705 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1190_l1158_DUPLICATE_9705_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_b856(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_4851_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_4851_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1190_l1158_DUPLICATE_9705_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l1190_l1158_DUPLICATE_9705_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
