-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity neq_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_226c8821;
architecture arch of neq_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1242_c6_2de8]
signal BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1242_c2_ba05]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1242_c2_ba05]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1242_c2_ba05]
signal result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1242_c2_ba05]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1242_c2_ba05]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1242_c2_ba05]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1242_c2_ba05]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1242_c2_ba05]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1242_c2_ba05]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1242_c2_ba05]
signal n8_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1242_c2_ba05]
signal t8_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1255_c11_4a49]
signal BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1255_c7_9645]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1255_c7_9645]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1255_c7_9645]
signal result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1255_c7_9645]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1255_c7_9645]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1255_c7_9645]
signal n8_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1255_c7_9645]
signal t8_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1258_c11_49a0]
signal BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1258_c7_af82]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1258_c7_af82]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1258_c7_af82]
signal result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1258_c7_af82]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1258_c7_af82]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1258_c7_af82]
signal n8_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1258_c7_af82]
signal t8_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1261_c11_12c3]
signal BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1261_c7_4296]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1261_c7_4296]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1261_c7_4296]
signal result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1261_c7_4296]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1261_c7_4296]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1261_c7_4296]
signal n8_MUX_uxn_opcodes_h_l1261_c7_4296_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1261_c7_4296_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1263_c30_ab4a]
signal sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1266_c21_470a]
signal BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1266_c21_eecb]
signal MUX_uxn_opcodes_h_l1266_c21_eecb_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1266_c21_eecb_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1266_c21_eecb_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1266_c21_eecb_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8
BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_left,
BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_right,
BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_cond,
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output);

-- n8_MUX_uxn_opcodes_h_l1242_c2_ba05
n8_MUX_uxn_opcodes_h_l1242_c2_ba05 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1242_c2_ba05_cond,
n8_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue,
n8_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse,
n8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output);

-- t8_MUX_uxn_opcodes_h_l1242_c2_ba05
t8_MUX_uxn_opcodes_h_l1242_c2_ba05 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1242_c2_ba05_cond,
t8_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue,
t8_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse,
t8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49
BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_left,
BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_right,
BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_cond,
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_return_output);

-- n8_MUX_uxn_opcodes_h_l1255_c7_9645
n8_MUX_uxn_opcodes_h_l1255_c7_9645 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1255_c7_9645_cond,
n8_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue,
n8_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse,
n8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output);

-- t8_MUX_uxn_opcodes_h_l1255_c7_9645
t8_MUX_uxn_opcodes_h_l1255_c7_9645 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1255_c7_9645_cond,
t8_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue,
t8_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse,
t8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0
BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_left,
BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_right,
BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_cond,
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_return_output);

-- n8_MUX_uxn_opcodes_h_l1258_c7_af82
n8_MUX_uxn_opcodes_h_l1258_c7_af82 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1258_c7_af82_cond,
n8_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue,
n8_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse,
n8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output);

-- t8_MUX_uxn_opcodes_h_l1258_c7_af82
t8_MUX_uxn_opcodes_h_l1258_c7_af82 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1258_c7_af82_cond,
t8_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue,
t8_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse,
t8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3
BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_left,
BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_right,
BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_cond,
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_return_output);

-- n8_MUX_uxn_opcodes_h_l1261_c7_4296
n8_MUX_uxn_opcodes_h_l1261_c7_4296 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1261_c7_4296_cond,
n8_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue,
n8_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse,
n8_MUX_uxn_opcodes_h_l1261_c7_4296_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a
sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_ins,
sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_x,
sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_y,
sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a
BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_left,
BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_right,
BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_return_output);

-- MUX_uxn_opcodes_h_l1266_c21_eecb
MUX_uxn_opcodes_h_l1266_c21_eecb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1266_c21_eecb_cond,
MUX_uxn_opcodes_h_l1266_c21_eecb_iftrue,
MUX_uxn_opcodes_h_l1266_c21_eecb_iffalse,
MUX_uxn_opcodes_h_l1266_c21_eecb_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
 n8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
 t8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_return_output,
 n8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output,
 t8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_return_output,
 n8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output,
 t8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_return_output,
 n8_MUX_uxn_opcodes_h_l1261_c7_4296_return_output,
 sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_return_output,
 MUX_uxn_opcodes_h_l1266_c21_eecb_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1247_c3_8a14 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1252_c3_d7bd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1242_c2_ba05_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1256_c3_9b61 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1255_c7_9645_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1261_c7_4296_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1258_c7_af82_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1265_c3_9f90 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1261_c7_4296_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1266_c21_eecb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1266_c21_eecb_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1266_c21_eecb_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1266_c21_eecb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_cf00_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_a9b6_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_d87d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_79f5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_0393_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1238_l1270_DUPLICATE_0ec7_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1252_c3_d7bd := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1252_c3_d7bd;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1265_c3_9f90 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1265_c3_9f90;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1266_c21_eecb_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_MUX_uxn_opcodes_h_l1266_c21_eecb_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1256_c3_9b61 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1256_c3_9b61;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1247_c3_8a14 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1247_c3_8a14;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_a9b6 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_a9b6_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_cf00 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_cf00_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_79f5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_79f5_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1261_c11_12c3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1242_c2_ba05_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1242_c6_2de8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1266_c21_470a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1242_c2_ba05_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_0393 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_0393_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1255_c11_4a49] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_left;
     BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_return_output := BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1258_c11_49a0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1242_c2_ba05_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_d87d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_d87d_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l1263_c30_ab4a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_ins;
     sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_x;
     sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_return_output := sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1242_c2_ba05_return_output := result.is_stack_index_flipped;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1242_c2_ba05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1242_c2_ba05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_2de8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1255_c7_9645_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1255_c7_9645_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_4a49_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1258_c7_af82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1258_c7_af82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_49a0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1261_c7_4296_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_12c3_return_output;
     VAR_MUX_uxn_opcodes_h_l1266_c21_eecb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_470a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_a9b6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_a9b6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_a9b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_79f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_79f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_79f5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_d87d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_d87d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_d87d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_0393_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_0393_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_cf00_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_cf00_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_cf00_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_cf00_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1242_c2_ba05_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1242_c2_ba05_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1242_c2_ba05_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1242_c2_ba05_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_ab4a_return_output;
     -- t8_MUX[uxn_opcodes_h_l1258_c7_af82] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1258_c7_af82_cond <= VAR_t8_MUX_uxn_opcodes_h_l1258_c7_af82_cond;
     t8_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue;
     t8_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output := t8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1261_c7_4296] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_return_output;

     -- n8_MUX[uxn_opcodes_h_l1261_c7_4296] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1261_c7_4296_cond <= VAR_n8_MUX_uxn_opcodes_h_l1261_c7_4296_cond;
     n8_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue;
     n8_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1261_c7_4296_return_output := n8_MUX_uxn_opcodes_h_l1261_c7_4296_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1261_c7_4296] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1261_c7_4296] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_return_output;

     -- MUX[uxn_opcodes_h_l1266_c21_eecb] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1266_c21_eecb_cond <= VAR_MUX_uxn_opcodes_h_l1266_c21_eecb_cond;
     MUX_uxn_opcodes_h_l1266_c21_eecb_iftrue <= VAR_MUX_uxn_opcodes_h_l1266_c21_eecb_iftrue;
     MUX_uxn_opcodes_h_l1266_c21_eecb_iffalse <= VAR_MUX_uxn_opcodes_h_l1266_c21_eecb_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1266_c21_eecb_return_output := MUX_uxn_opcodes_h_l1266_c21_eecb_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1261_c7_4296] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue := VAR_MUX_uxn_opcodes_h_l1266_c21_eecb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1261_c7_4296_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_4296_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_4296_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_4296_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_4296_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1258_c7_af82] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1258_c7_af82] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;

     -- n8_MUX[uxn_opcodes_h_l1258_c7_af82] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1258_c7_af82_cond <= VAR_n8_MUX_uxn_opcodes_h_l1258_c7_af82_cond;
     n8_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue;
     n8_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output := n8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;

     -- t8_MUX[uxn_opcodes_h_l1255_c7_9645] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1255_c7_9645_cond <= VAR_t8_MUX_uxn_opcodes_h_l1255_c7_9645_cond;
     t8_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue;
     t8_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output := t8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1258_c7_af82] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1258_c7_af82] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1261_c7_4296] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_return_output := result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_4296_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1255_c7_9645] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1255_c7_9645] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1255_c7_9645] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1255_c7_9645] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;

     -- n8_MUX[uxn_opcodes_h_l1255_c7_9645] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1255_c7_9645_cond <= VAR_n8_MUX_uxn_opcodes_h_l1255_c7_9645_cond;
     n8_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue;
     n8_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output := n8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;

     -- t8_MUX[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1242_c2_ba05_cond <= VAR_t8_MUX_uxn_opcodes_h_l1242_c2_ba05_cond;
     t8_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue;
     t8_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output := t8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1258_c7_af82] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_return_output := result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_af82_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output;
     -- n8_MUX[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1242_c2_ba05_cond <= VAR_n8_MUX_uxn_opcodes_h_l1242_c2_ba05_cond;
     n8_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue;
     n8_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output := n8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1255_c7_9645] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_return_output := result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_9645_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1242_c2_ba05] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output := result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1238_l1270_DUPLICATE_0ec7 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1238_l1270_DUPLICATE_0ec7_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_ba05_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1238_l1270_DUPLICATE_0ec7_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1238_l1270_DUPLICATE_0ec7_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
