-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity opc_sub_phased_0CLK_c3dfc98c is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_sub_phased_0CLK_c3dfc98c;
architecture arch of opc_sub_phased_0CLK_c3dfc98c is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l1041_c6_9b00]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1041_c1_4dd3]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1044_c7_5385]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1041_c2_74e2]
signal t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1041_c2_74e2]
signal n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1041_c2_74e2]
signal result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output : unsigned(0 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l1042_c12_dd02]
signal set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1044_c11_a9df]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1044_c1_821b]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1047_c7_0d7f]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1044_c7_5385]
signal t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1044_c7_5385]
signal n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1044_c7_5385]
signal result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output : unsigned(0 downto 0);

-- t_register[uxn_opcodes_phased_h_l1045_c8_bc21]
signal t_register_uxn_opcodes_phased_h_l1045_c8_bc21_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l1045_c8_bc21_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l1045_c8_bc21_stack_ptr : unsigned(7 downto 0);
signal t_register_uxn_opcodes_phased_h_l1045_c8_bc21_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1047_c11_4e93]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1047_c1_3388]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1050_c7_5743]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1047_c7_0d7f]
signal t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1047_c7_0d7f]
signal n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1047_c7_0d7f]
signal result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l1048_c8_4d61]
signal n_register_uxn_opcodes_phased_h_l1048_c8_4d61_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1048_c8_4d61_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1048_c8_4d61_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l1048_c8_4d61_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1050_c11_a996]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1050_c1_8d64]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1053_c7_7a8a]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1050_c7_5743]
signal n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1050_c7_5743]
signal result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l1051_c8_634c]
signal n_register_uxn_opcodes_phased_h_l1051_c8_634c_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1051_c8_634c_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1051_c8_634c_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l1051_c8_634c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1053_c11_96c7]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1053_c1_c123]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1056_c7_04d1]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1053_c7_7a8a]
signal result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output : unsigned(0 downto 0);

-- set[uxn_opcodes_phased_h_l1054_c3_837c]
signal set_uxn_opcodes_phased_h_l1054_c3_837c_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l1054_c3_837c_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1054_c3_837c_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l1054_c3_837c_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1054_c3_837c_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1054_c3_837c_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1054_c3_837c_add : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1056_c11_3187]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1056_c1_0e0e]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1056_c7_04d1]
signal result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output : unsigned(0 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_phased_h_l1057_c33_4fa0]
signal BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_return_output : unsigned(7 downto 0);

-- put_stack[uxn_opcodes_phased_h_l1057_c3_8590]
signal put_stack_uxn_opcodes_phased_h_l1057_c3_8590_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1057_c3_8590_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1057_c3_8590_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1057_c3_8590_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1057_c3_8590_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1059_c11_16b2]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1059_c7_455e]
signal result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00
BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2
t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond,
t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2
n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond,
n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2
result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond,
result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue,
result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse,
result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02
set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02 : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_sp,
set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_k,
set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_mul,
set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_add,
set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df
BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385
t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond,
t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385
n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond,
n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1044_c7_5385
result_MUX_uxn_opcodes_phased_h_l1044_c7_5385 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond,
result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue,
result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse,
result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output);

-- t_register_uxn_opcodes_phased_h_l1045_c8_bc21
t_register_uxn_opcodes_phased_h_l1045_c8_bc21 : entity work.t_register_0CLK_621d5f60 port map (
clk,
t_register_uxn_opcodes_phased_h_l1045_c8_bc21_CLOCK_ENABLE,
t_register_uxn_opcodes_phased_h_l1045_c8_bc21_stack_index,
t_register_uxn_opcodes_phased_h_l1045_c8_bc21_stack_ptr,
t_register_uxn_opcodes_phased_h_l1045_c8_bc21_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93
BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f
t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond,
t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f
n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond,
n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f
result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond,
result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue,
result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse,
result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output);

-- n_register_uxn_opcodes_phased_h_l1048_c8_4d61
n_register_uxn_opcodes_phased_h_l1048_c8_4d61 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l1048_c8_4d61_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l1048_c8_4d61_stack_index,
n_register_uxn_opcodes_phased_h_l1048_c8_4d61_stack_ptr,
n_register_uxn_opcodes_phased_h_l1048_c8_4d61_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996
BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743
n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond,
n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1050_c7_5743
result_MUX_uxn_opcodes_phased_h_l1050_c7_5743 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond,
result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue,
result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse,
result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output);

-- n_register_uxn_opcodes_phased_h_l1051_c8_634c
n_register_uxn_opcodes_phased_h_l1051_c8_634c : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l1051_c8_634c_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l1051_c8_634c_stack_index,
n_register_uxn_opcodes_phased_h_l1051_c8_634c_stack_ptr,
n_register_uxn_opcodes_phased_h_l1051_c8_634c_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7
BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a
result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_cond,
result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iftrue,
result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iffalse,
result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output);

-- set_uxn_opcodes_phased_h_l1054_c3_837c
set_uxn_opcodes_phased_h_l1054_c3_837c : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l1054_c3_837c_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l1054_c3_837c_sp,
set_uxn_opcodes_phased_h_l1054_c3_837c_stack_index,
set_uxn_opcodes_phased_h_l1054_c3_837c_ins,
set_uxn_opcodes_phased_h_l1054_c3_837c_k,
set_uxn_opcodes_phased_h_l1054_c3_837c_mul,
set_uxn_opcodes_phased_h_l1054_c3_837c_add);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187
BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1
result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_cond,
result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iftrue,
result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iffalse,
result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output);

-- BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0
BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_left,
BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_right,
BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_return_output);

-- put_stack_uxn_opcodes_phased_h_l1057_c3_8590
put_stack_uxn_opcodes_phased_h_l1057_c3_8590 : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l1057_c3_8590_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l1057_c3_8590_sp,
put_stack_uxn_opcodes_phased_h_l1057_c3_8590_stack_index,
put_stack_uxn_opcodes_phased_h_l1057_c3_8590_offset,
put_stack_uxn_opcodes_phased_h_l1057_c3_8590_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2
BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1059_c7_455e
result_MUX_uxn_opcodes_phased_h_l1059_c7_455e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_cond,
result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_iftrue,
result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_iffalse,
result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 n8,
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output,
 result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output,
 set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output,
 result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output,
 t_register_uxn_opcodes_phased_h_l1045_c8_bc21_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output,
 result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output,
 n_register_uxn_opcodes_phased_h_l1048_c8_4d61_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output,
 result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output,
 n_register_uxn_opcodes_phased_h_l1051_c8_634c_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output,
 result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_return_output,
 result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output,
 BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_return_output,
 result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1045_c8_bc21_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1045_c8_bc21_stack_ptr : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1045_c8_bc21_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1045_c8_bc21_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1048_c8_4d61_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1048_c8_4d61_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1048_c8_4d61_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1048_c8_4d61_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1051_c8_634c_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1051_c8_634c_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1051_c8_634c_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1051_c8_634c_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_cond : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_value : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_return_output : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_n8 := n8;
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_mul := resize(to_unsigned(2, 2), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_right := to_unsigned(5, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue := to_unsigned(0, 1);
     VAR_result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_right := to_unsigned(1, 1);
     VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_offset := resize(to_unsigned(0, 1), 8);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_right := to_unsigned(6, 3);
     VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_add := resize(to_signed(-1, 2), 8);
     VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_add := resize(to_signed(-1, 2), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_right := to_unsigned(2, 2);
     VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_mul := resize(to_unsigned(2, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_k := VAR_k;
     VAR_BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_left := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_left := VAR_phase;
     VAR_result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_iffalse := result;
     VAR_n_register_uxn_opcodes_phased_h_l1048_c8_4d61_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l1051_c8_634c_stack_ptr := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_sp := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_sp := VAR_sp;
     VAR_t_register_uxn_opcodes_phased_h_l1045_c8_bc21_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l1048_c8_4d61_stack_index := VAR_stack_index;
     VAR_n_register_uxn_opcodes_phased_h_l1051_c8_634c_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_phased_h_l1045_c8_bc21_stack_index := VAR_stack_index;
     VAR_BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_right := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1050_c11_a996] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1056_c11_3187] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1053_c11_96c7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1044_c11_a9df] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1041_c6_9b00] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_return_output;

     -- BIN_OP_MINUS[uxn_opcodes_phased_h_l1057_c33_4fa0] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_left <= VAR_BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_left;
     BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_right <= VAR_BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_return_output := BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1047_c11_4e93] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1059_c11_16b2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1041_c6_9b00_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1044_c11_a9df_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1047_c11_4e93_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1050_c11_a996_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1053_c11_96c7_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1056_c11_3187_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1059_c11_16b2_return_output;
     VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_value := VAR_BIN_OP_MINUS_uxn_opcodes_phased_h_l1057_c33_4fa0_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l1059_c7_455e] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_cond;
     result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_return_output := result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1044_c7_5385] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1041_c1_4dd3] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1041_c1_4dd3_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1059_c7_455e_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l1056_c7_04d1] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_cond;
     result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output := result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1047_c7_0d7f] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output;

     -- set_will_fail[uxn_opcodes_phased_h_l1042_c12_dd02] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_sp;
     set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_k;
     set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_mul;
     set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_return_output := set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1044_c1_821b] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output;
     VAR_t_register_uxn_opcodes_phased_h_l1045_c8_bc21_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1044_c1_821b_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l1042_c12_dd02_return_output;
     -- t_register[uxn_opcodes_phased_h_l1045_c8_bc21] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_phased_h_l1045_c8_bc21_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_phased_h_l1045_c8_bc21_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_phased_h_l1045_c8_bc21_stack_index <= VAR_t_register_uxn_opcodes_phased_h_l1045_c8_bc21_stack_index;
     t_register_uxn_opcodes_phased_h_l1045_c8_bc21_stack_ptr <= VAR_t_register_uxn_opcodes_phased_h_l1045_c8_bc21_stack_ptr;
     -- Outputs
     VAR_t_register_uxn_opcodes_phased_h_l1045_c8_bc21_return_output := t_register_uxn_opcodes_phased_h_l1045_c8_bc21_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1053_c7_7a8a] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_cond;
     result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output := result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1047_c1_3388] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1050_c7_5743] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l1048_c8_4d61_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1047_c1_3388_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue := VAR_t_register_uxn_opcodes_phased_h_l1045_c8_bc21_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1050_c1_8d64] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1050_c7_5743] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond;
     result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output := result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1053_c7_7a8a] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output;

     -- n_register[uxn_opcodes_phased_h_l1048_c8_4d61] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l1048_c8_4d61_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l1048_c8_4d61_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l1048_c8_4d61_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l1048_c8_4d61_stack_index;
     n_register_uxn_opcodes_phased_h_l1048_c8_4d61_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l1048_c8_4d61_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l1048_c8_4d61_return_output := n_register_uxn_opcodes_phased_h_l1048_c8_4d61_return_output;

     -- Submodule level 5
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c7_7a8a_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l1051_c8_634c_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1050_c1_8d64_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue := VAR_n_register_uxn_opcodes_phased_h_l1048_c8_4d61_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output;
     -- t8_MUX[uxn_opcodes_phased_h_l1047_c7_0d7f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond;
     t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output := t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1056_c7_04d1] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output;

     -- n_register[uxn_opcodes_phased_h_l1051_c8_634c] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l1051_c8_634c_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l1051_c8_634c_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l1051_c8_634c_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l1051_c8_634c_stack_index;
     n_register_uxn_opcodes_phased_h_l1051_c8_634c_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l1051_c8_634c_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l1051_c8_634c_return_output := n_register_uxn_opcodes_phased_h_l1051_c8_634c_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1047_c7_0d7f] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond;
     result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output := result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1053_c1_c123] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_return_output;

     -- Submodule level 6
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c7_04d1_return_output;
     VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1053_c1_c123_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue := VAR_n_register_uxn_opcodes_phased_h_l1051_c8_634c_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1050_c7_5743] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_cond;
     n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output := n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output;

     -- set[uxn_opcodes_phased_h_l1054_c3_837c] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l1054_c3_837c_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l1054_c3_837c_sp <= VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_sp;
     set_uxn_opcodes_phased_h_l1054_c3_837c_stack_index <= VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_stack_index;
     set_uxn_opcodes_phased_h_l1054_c3_837c_ins <= VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_ins;
     set_uxn_opcodes_phased_h_l1054_c3_837c_k <= VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_k;
     set_uxn_opcodes_phased_h_l1054_c3_837c_mul <= VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_mul;
     set_uxn_opcodes_phased_h_l1054_c3_837c_add <= VAR_set_uxn_opcodes_phased_h_l1054_c3_837c_add;
     -- Outputs

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1056_c1_0e0e] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l1044_c7_5385] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond;
     t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output := t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1044_c7_5385] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond;
     result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output := result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output;

     -- Submodule level 7
     VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1056_c1_0e0e_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1050_c7_5743_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1047_c7_0d7f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_cond;
     n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output := n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output;

     -- put_stack[uxn_opcodes_phased_h_l1057_c3_8590] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l1057_c3_8590_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l1057_c3_8590_sp <= VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_sp;
     put_stack_uxn_opcodes_phased_h_l1057_c3_8590_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_stack_index;
     put_stack_uxn_opcodes_phased_h_l1057_c3_8590_offset <= VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_offset;
     put_stack_uxn_opcodes_phased_h_l1057_c3_8590_value <= VAR_put_stack_uxn_opcodes_phased_h_l1057_c3_8590_value;
     -- Outputs

     -- result_MUX[uxn_opcodes_phased_h_l1041_c2_74e2] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond;
     result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output := result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l1041_c2_74e2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond;
     t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output := t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output;

     -- Submodule level 8
     VAR_n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1047_c7_0d7f_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1044_c7_5385] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_cond;
     n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output := n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output;

     -- Submodule level 9
     VAR_n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1044_c7_5385_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1041_c2_74e2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_cond;
     n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output := n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output;

     -- Submodule level 10
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_phased_h_l1041_c2_74e2_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     n8 <= REG_COMB_n8;
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
