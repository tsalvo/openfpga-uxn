-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 56
entity inc2_0CLK_a6885b22 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc2_0CLK_a6885b22;
architecture arch of inc2_0CLK_a6885b22 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1291_c6_8fe5]
signal BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1291_c1_eeca]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1291_c2_d9cb]
signal tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1291_c2_d9cb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1291_c2_d9cb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1291_c2_d9cb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1291_c2_d9cb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1291_c2_d9cb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1291_c2_d9cb]
signal result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l1291_c2_d9cb]
signal t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l1292_c3_440e[uxn_opcodes_h_l1292_c3_440e]
signal printf_uxn_opcodes_h_l1292_c3_440e_uxn_opcodes_h_l1292_c3_440e_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1296_c11_1b4c]
signal BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1296_c7_314f]
signal tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1296_c7_314f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1296_c7_314f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1296_c7_314f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1296_c7_314f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1296_c7_314f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1296_c7_314f]
signal result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l1296_c7_314f]
signal t16_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1299_c11_a61f]
signal BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1299_c7_ad11]
signal tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1299_c7_ad11]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1299_c7_ad11]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1299_c7_ad11]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1299_c7_ad11]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1299_c7_ad11]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1299_c7_ad11]
signal result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l1299_c7_ad11]
signal t16_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l1301_c3_d0d4]
signal CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1303_c11_a708]
signal BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1303_c7_b859]
signal tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1303_c7_b859]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1303_c7_b859]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1303_c7_b859]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1303_c7_b859]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1303_c7_b859]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1303_c7_b859]
signal result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l1303_c7_b859]
signal t16_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l1304_c3_30f6]
signal BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1305_c11_7f9a]
signal BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_return_output : unsigned(16 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1307_c30_58a4]
signal sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1312_c11_2a17]
signal BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1312_c7_55c1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1312_c7_55c1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1312_c7_55c1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1312_c7_55c1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1312_c7_55c1]
signal result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output : unsigned(7 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l1315_c31_6921]
signal CONST_SR_8_uxn_opcodes_h_l1315_c31_6921_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l1315_c31_6921_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1317_c11_b740]
signal BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1317_c7_1093]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1317_c7_1093]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_4e73( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5
BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_left,
BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_right,
BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb
tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond,
tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue,
tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse,
tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb
result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb
result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb
result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb
result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb
result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond,
result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output);

-- t16_MUX_uxn_opcodes_h_l1291_c2_d9cb
t16_MUX_uxn_opcodes_h_l1291_c2_d9cb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond,
t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue,
t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse,
t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output);

-- printf_uxn_opcodes_h_l1292_c3_440e_uxn_opcodes_h_l1292_c3_440e
printf_uxn_opcodes_h_l1292_c3_440e_uxn_opcodes_h_l1292_c3_440e : entity work.printf_uxn_opcodes_h_l1292_c3_440e_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1292_c3_440e_uxn_opcodes_h_l1292_c3_440e_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c
BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_left,
BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_right,
BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1296_c7_314f
tmp16_MUX_uxn_opcodes_h_l1296_c7_314f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_cond,
tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue,
tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse,
tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f
result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f
result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f
result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f
result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_return_output);

-- t16_MUX_uxn_opcodes_h_l1296_c7_314f
t16_MUX_uxn_opcodes_h_l1296_c7_314f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1296_c7_314f_cond,
t16_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue,
t16_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse,
t16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f
BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_left,
BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_right,
BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11
tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_cond,
tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue,
tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse,
tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11
result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11
result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_cond,
result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output);

-- t16_MUX_uxn_opcodes_h_l1299_c7_ad11
t16_MUX_uxn_opcodes_h_l1299_c7_ad11 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1299_c7_ad11_cond,
t16_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue,
t16_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse,
t16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output);

-- CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4
CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4_x,
CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708
BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_left,
BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_right,
BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1303_c7_b859
tmp16_MUX_uxn_opcodes_h_l1303_c7_b859 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_cond,
tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue,
tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse,
tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859
result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859
result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859
result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859
result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859
result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_cond,
result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_return_output);

-- t16_MUX_uxn_opcodes_h_l1303_c7_b859
t16_MUX_uxn_opcodes_h_l1303_c7_b859 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1303_c7_b859_cond,
t16_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue,
t16_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse,
t16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6
BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_left,
BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_right,
BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a
BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_left,
BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_right,
BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4
sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_ins,
sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_x,
sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_y,
sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17
BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_left,
BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_right,
BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1
result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1
result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1
result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1
result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_cond,
result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output);

-- CONST_SR_8_uxn_opcodes_h_l1315_c31_6921
CONST_SR_8_uxn_opcodes_h_l1315_c31_6921 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l1315_c31_6921_x,
CONST_SR_8_uxn_opcodes_h_l1315_c31_6921_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740
BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_left,
BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_right,
BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_return_output,
 tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output,
 t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output,
 tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_return_output,
 t16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output,
 tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output,
 t16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output,
 CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output,
 tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_return_output,
 t16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output,
 BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_return_output,
 sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output,
 CONST_SR_8_uxn_opcodes_h_l1315_c31_6921_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_iffalse : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1293_c3_a4f1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1292_c3_440e_uxn_opcodes_h_l1292_c3_440e_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1297_c3_efed : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1296_c7_314f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1299_c7_ad11_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_uxn_opcodes_h_l1305_c3_53d5 : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1309_c3_e63e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1303_c7_b859_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_return_output : unsigned(16 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1310_c21_fda8_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1314_c3_7641 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l1315_c31_6921_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l1315_c31_6921_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1315_c21_6997_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1312_l1299_l1296_l1291_DUPLICATE_a4ec_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_96c1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1299_l1291_l1303_l1296_DUPLICATE_91aa_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_be15_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1317_l1312_l1303_l1299_l1296_DUPLICATE_560a_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1304_l1300_DUPLICATE_b59e_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1299_l1312_DUPLICATE_95b5_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1287_l1322_DUPLICATE_06ea_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1297_c3_efed := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1297_c3_efed;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_iffalse := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1314_c3_7641 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1314_c3_7641;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1309_c3_e63e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1309_c3_e63e;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1293_c3_a4f1 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1293_c3_a4f1;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse := t16;
     VAR_CONST_SR_8_uxn_opcodes_h_l1315_c31_6921_x := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse := tmp16;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1299_l1291_l1303_l1296_DUPLICATE_91aa LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1299_l1291_l1303_l1296_DUPLICATE_91aa_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1312_l1299_l1296_l1291_DUPLICATE_a4ec LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1312_l1299_l1296_l1291_DUPLICATE_a4ec_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l1307_c30_58a4] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_ins;
     sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_x;
     sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_return_output := sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1312_c11_2a17] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_left;
     BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_return_output := BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_be15 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_be15_return_output := result.u8_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1299_l1312_DUPLICATE_95b5 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1299_l1312_DUPLICATE_95b5_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1303_c11_a708] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_left;
     BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output := BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1317_c11_b740] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_left;
     BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_return_output := BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_return_output;

     -- CONST_SR_8[uxn_opcodes_h_l1315_c31_6921] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l1315_c31_6921_x <= VAR_CONST_SR_8_uxn_opcodes_h_l1315_c31_6921_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l1315_c31_6921_return_output := CONST_SR_8_uxn_opcodes_h_l1315_c31_6921_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_96c1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_96c1_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1291_c6_8fe5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1299_c11_a61f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1317_l1312_l1303_l1299_l1296_DUPLICATE_560a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1317_l1312_l1303_l1299_l1296_DUPLICATE_560a_return_output := result.is_opc_done;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1304_l1300_DUPLICATE_b59e LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1304_l1300_DUPLICATE_b59e_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1296_c11_1b4c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_8fe5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1296_c7_314f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_1b4c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1299_c7_ad11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_a61f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1303_c7_b859_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_a708_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_2a17_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_b740_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1304_l1300_DUPLICATE_b59e_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1304_l1300_DUPLICATE_b59e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1299_l1291_l1303_l1296_DUPLICATE_91aa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1299_l1291_l1303_l1296_DUPLICATE_91aa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1299_l1291_l1303_l1296_DUPLICATE_91aa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1299_l1291_l1303_l1296_DUPLICATE_91aa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1317_l1312_l1303_l1299_l1296_DUPLICATE_560a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1317_l1312_l1303_l1299_l1296_DUPLICATE_560a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1317_l1312_l1303_l1299_l1296_DUPLICATE_560a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1317_l1312_l1303_l1299_l1296_DUPLICATE_560a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1317_l1312_l1303_l1299_l1296_DUPLICATE_560a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_96c1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_96c1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_96c1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_96c1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1312_l1299_l1296_l1291_DUPLICATE_a4ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1312_l1299_l1296_l1291_DUPLICATE_a4ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1312_l1299_l1296_l1291_DUPLICATE_a4ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1312_l1299_l1296_l1291_DUPLICATE_a4ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1312_l1299_l1296_l1291_DUPLICATE_a4ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1299_l1312_DUPLICATE_95b5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1299_l1312_DUPLICATE_95b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_be15_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_be15_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_be15_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1299_l1291_l1296_l1312_DUPLICATE_be15_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_58a4_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1317_c7_1093] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1312_c7_55c1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1312_c7_55c1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l1315_c21_6997] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1315_c21_6997_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l1315_c31_6921_return_output);

     -- CONST_SL_8[uxn_opcodes_h_l1301_c3_d0d4] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4_x <= VAR_CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4_return_output := CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1291_c1_eeca] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l1304_c3_30f6] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_left;
     BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_return_output := BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1317_c7_1093] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1303_c7_b859] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;

     -- Submodule level 2
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_left := VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_30f6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1315_c21_6997_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l1301_c3_d0d4_return_output;
     VAR_printf_uxn_opcodes_h_l1292_c3_440e_uxn_opcodes_h_l1292_c3_440e_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_eeca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_1093_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_1093_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output;
     -- t16_MUX[uxn_opcodes_h_l1303_c7_b859] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1303_c7_b859_cond <= VAR_t16_MUX_uxn_opcodes_h_l1303_c7_b859_cond;
     t16_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue;
     t16_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output := t16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1305_c11_7f9a] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_return_output;

     -- printf_uxn_opcodes_h_l1292_c3_440e[uxn_opcodes_h_l1292_c3_440e] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1292_c3_440e_uxn_opcodes_h_l1292_c3_440e_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1292_c3_440e_uxn_opcodes_h_l1292_c3_440e_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1299_c7_ad11] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1303_c7_b859] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1312_c7_55c1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1312_c7_55c1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1303_c7_b859] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1312_c7_55c1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output := result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output;

     -- Submodule level 3
     VAR_tmp16_uxn_opcodes_h_l1305_c3_53d5 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_7f9a_return_output, 16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_55c1_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue := VAR_tmp16_uxn_opcodes_h_l1305_c3_53d5;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1299_c7_ad11] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1303_c7_b859] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1303_c7_b859] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1299_c7_ad11] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l1310_c21_fda8] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1310_c21_fda8_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_tmp16_uxn_opcodes_h_l1305_c3_53d5);

     -- t16_MUX[uxn_opcodes_h_l1299_c7_ad11] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1299_c7_ad11_cond <= VAR_t16_MUX_uxn_opcodes_h_l1299_c7_ad11_cond;
     t16_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue;
     t16_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output := t16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1303_c7_b859] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_cond;
     tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output := tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1296_c7_314f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;

     -- Submodule level 4
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1310_c21_fda8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;
     -- t16_MUX[uxn_opcodes_h_l1296_c7_314f] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1296_c7_314f_cond <= VAR_t16_MUX_uxn_opcodes_h_l1296_c7_314f_cond;
     t16_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue;
     t16_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output := t16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1303_c7_b859] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_return_output := result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1299_c7_ad11] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1296_c7_314f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1291_c2_d9cb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1299_c7_ad11] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_cond;
     tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output := tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1299_c7_ad11] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1296_c7_314f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_b859_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1296_c7_314f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1296_c7_314f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1291_c2_d9cb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1291_c2_d9cb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output;

     -- t16_MUX[uxn_opcodes_h_l1291_c2_d9cb] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond <= VAR_t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond;
     t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue;
     t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output := t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1296_c7_314f] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_cond;
     tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output := tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1299_c7_ad11] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output := result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_ad11_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1291_c2_d9cb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1291_c2_d9cb] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond;
     tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output := tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1291_c2_d9cb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1296_c7_314f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;

     -- Submodule level 7
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_314f_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1291_c2_d9cb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output := result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1287_l1322_DUPLICATE_06ea LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1287_l1322_DUPLICATE_06ea_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4e73(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_d9cb_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1287_l1322_DUPLICATE_06ea_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1287_l1322_DUPLICATE_06ea_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
