-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 49
entity ora2_0CLK_06b39b76 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end ora2_0CLK_06b39b76;
architecture arch of ora2_0CLK_06b39b76 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l953_c6_0b67]
signal BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l953_c2_af81]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l953_c2_af81]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l953_c2_af81]
signal result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l953_c2_af81]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l953_c2_af81]
signal result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l953_c2_af81]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l953_c2_af81]
signal result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l953_c2_af81]
signal n16_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l953_c2_af81]
signal tmp16_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l953_c2_af81]
signal t16_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l961_c11_bb22]
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l961_c7_0f37]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l961_c7_0f37]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l961_c7_0f37]
signal result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l961_c7_0f37]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l961_c7_0f37]
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l961_c7_0f37]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l961_c7_0f37]
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l961_c7_0f37]
signal n16_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l961_c7_0f37]
signal tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l961_c7_0f37]
signal t16_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l964_c11_42ac]
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l964_c7_0bed]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l964_c7_0bed]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l964_c7_0bed]
signal result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l964_c7_0bed]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l964_c7_0bed]
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l964_c7_0bed]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l964_c7_0bed]
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l964_c7_0bed]
signal n16_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l964_c7_0bed]
signal tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l964_c7_0bed]
signal t16_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l967_c30_2d64]
signal sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l969_c11_6204]
signal BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l969_c7_8db1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l969_c7_8db1]
signal result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l969_c7_8db1]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l969_c7_8db1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l969_c7_8db1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l969_c7_8db1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l969_c7_8db1]
signal n16_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l969_c7_8db1]
signal tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l971_c11_a04b]
signal BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l977_c11_6816]
signal BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l977_c7_bbfe]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l977_c7_bbfe]
signal result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l977_c7_bbfe]
signal result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67
BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_left,
BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_right,
BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81
result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81
result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_cond,
result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81
result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81
result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81
result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_return_output);

-- n16_MUX_uxn_opcodes_h_l953_c2_af81
n16_MUX_uxn_opcodes_h_l953_c2_af81 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l953_c2_af81_cond,
n16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue,
n16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse,
n16_MUX_uxn_opcodes_h_l953_c2_af81_return_output);

-- tmp16_MUX_uxn_opcodes_h_l953_c2_af81
tmp16_MUX_uxn_opcodes_h_l953_c2_af81 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l953_c2_af81_cond,
tmp16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue,
tmp16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse,
tmp16_MUX_uxn_opcodes_h_l953_c2_af81_return_output);

-- t16_MUX_uxn_opcodes_h_l953_c2_af81
t16_MUX_uxn_opcodes_h_l953_c2_af81 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l953_c2_af81_cond,
t16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue,
t16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse,
t16_MUX_uxn_opcodes_h_l953_c2_af81_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22
BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_left,
BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_right,
BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37
result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_cond,
result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_return_output);

-- n16_MUX_uxn_opcodes_h_l961_c7_0f37
n16_MUX_uxn_opcodes_h_l961_c7_0f37 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l961_c7_0f37_cond,
n16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue,
n16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse,
n16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output);

-- tmp16_MUX_uxn_opcodes_h_l961_c7_0f37
tmp16_MUX_uxn_opcodes_h_l961_c7_0f37 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_cond,
tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue,
tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse,
tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output);

-- t16_MUX_uxn_opcodes_h_l961_c7_0f37
t16_MUX_uxn_opcodes_h_l961_c7_0f37 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l961_c7_0f37_cond,
t16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue,
t16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse,
t16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac
BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_left,
BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_right,
BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed
result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_cond,
result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_return_output);

-- n16_MUX_uxn_opcodes_h_l964_c7_0bed
n16_MUX_uxn_opcodes_h_l964_c7_0bed : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l964_c7_0bed_cond,
n16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue,
n16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse,
n16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output);

-- tmp16_MUX_uxn_opcodes_h_l964_c7_0bed
tmp16_MUX_uxn_opcodes_h_l964_c7_0bed : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_cond,
tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue,
tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse,
tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output);

-- t16_MUX_uxn_opcodes_h_l964_c7_0bed
t16_MUX_uxn_opcodes_h_l964_c7_0bed : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l964_c7_0bed_cond,
t16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue,
t16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse,
t16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output);

-- sp_relative_shift_uxn_opcodes_h_l967_c30_2d64
sp_relative_shift_uxn_opcodes_h_l967_c30_2d64 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_ins,
sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_x,
sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_y,
sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204
BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_left,
BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_right,
BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1
result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1
result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_cond,
result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1
result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1
result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_return_output);

-- n16_MUX_uxn_opcodes_h_l969_c7_8db1
n16_MUX_uxn_opcodes_h_l969_c7_8db1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l969_c7_8db1_cond,
n16_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue,
n16_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse,
n16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output);

-- tmp16_MUX_uxn_opcodes_h_l969_c7_8db1
tmp16_MUX_uxn_opcodes_h_l969_c7_8db1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_cond,
tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue,
tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse,
tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b
BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_left,
BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_right,
BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816
BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_left,
BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_right,
BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe
result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe
result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
 n16_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
 tmp16_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
 t16_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_return_output,
 n16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output,
 tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output,
 t16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_return_output,
 n16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output,
 tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output,
 t16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output,
 sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_return_output,
 n16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output,
 tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output,
 BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_b59f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l953_c2_af81_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l953_c2_af81_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_d118 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l961_c7_0f37_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l964_c7_0bed_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l974_c3_8499 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l961_l953_l969_DUPLICATE_2a70_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l961_l964_l953_l969_DUPLICATE_92b8_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l961_l964_l953_DUPLICATE_e84b_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l977_l964_l953_DUPLICATE_0fc9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_6cef_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_c65d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l969_DUPLICATE_198d_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l983_l949_DUPLICATE_718c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_d118 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_d118;
     VAR_sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_y := resize(to_signed(-2, 3), 4);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_b59f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_b59f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l974_c3_8499 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l974_c3_8499;
     VAR_sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_right := to_unsigned(3, 2);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_left := VAR_previous_stack_read;
     VAR_n16_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_right := t16;
     VAR_t16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse := t16;
     VAR_tmp16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse := tmp16;
     -- BIN_OP_EQ[uxn_opcodes_h_l969_c11_6204] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_left;
     BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output := BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l977_c11_6816] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_left;
     BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_return_output := BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l961_l953_l969_DUPLICATE_2a70 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l961_l953_l969_DUPLICATE_2a70_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_c65d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_c65d_return_output := result.is_opc_done;

     -- BIN_OP_OR[uxn_opcodes_h_l971_c11_a04b] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_left;
     BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_return_output := BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l953_c6_0b67] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_left;
     BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output := BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l977_l964_l953_DUPLICATE_0fc9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l977_l964_l953_DUPLICATE_0fc9_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l961_c11_bb22] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_left;
     BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output := BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_6cef LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_6cef_return_output := result.is_stack_operation_16bit;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l961_l964_l953_DUPLICATE_e84b LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l961_l964_l953_DUPLICATE_e84b_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l961_l964_l953_l969_DUPLICATE_92b8 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l961_l964_l953_l969_DUPLICATE_92b8_return_output := result.u16_value;

     -- sp_relative_shift[uxn_opcodes_h_l967_c30_2d64] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_ins;
     sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_x <= VAR_sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_x;
     sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_y <= VAR_sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_return_output := sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l964_c11_42ac] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_left;
     BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output := BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l969_DUPLICATE_198d LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l969_DUPLICATE_198d_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_n16_MUX_uxn_opcodes_h_l953_c2_af81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l953_c2_af81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l953_c2_af81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c6_0b67_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l961_c7_0f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l961_c7_0f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_bb22_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l964_c7_0bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l964_c7_0bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_42ac_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l969_c7_8db1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l969_c11_6204_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l977_c11_6816_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l971_c11_a04b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l961_l964_l953_DUPLICATE_e84b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l961_l964_l953_DUPLICATE_e84b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l961_l964_l953_DUPLICATE_e84b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l961_l964_l953_l969_DUPLICATE_92b8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l961_l964_l953_l969_DUPLICATE_92b8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l961_l964_l953_l969_DUPLICATE_92b8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l961_l964_l953_l969_DUPLICATE_92b8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_c65d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_c65d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_c65d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_c65d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l961_l953_l969_DUPLICATE_2a70_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l961_l953_l969_DUPLICATE_2a70_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l961_l953_l969_DUPLICATE_2a70_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_6cef_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_6cef_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_6cef_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l961_l977_l964_l969_DUPLICATE_6cef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l977_l964_l953_DUPLICATE_0fc9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l977_l964_l953_DUPLICATE_0fc9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l977_l964_l953_DUPLICATE_0fc9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l977_l964_l953_DUPLICATE_0fc9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l969_DUPLICATE_198d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l969_DUPLICATE_198d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l967_c30_2d64_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l964_c7_0bed] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l969_c7_8db1] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_cond;
     tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue;
     tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output := tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l977_c7_bbfe] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l969_c7_8db1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l969_c7_8db1] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_cond;
     result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_return_output := result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l977_c7_bbfe] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output;

     -- n16_MUX[uxn_opcodes_h_l969_c7_8db1] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l969_c7_8db1_cond <= VAR_n16_MUX_uxn_opcodes_h_l969_c7_8db1_cond;
     n16_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue;
     n16_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output := n16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;

     -- t16_MUX[uxn_opcodes_h_l964_c7_0bed] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l964_c7_0bed_cond <= VAR_t16_MUX_uxn_opcodes_h_l964_c7_0bed_cond;
     t16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue;
     t16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output := t16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l969_c7_8db1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l977_c7_bbfe] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output;

     -- Submodule level 2
     VAR_n16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse := VAR_n16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l977_c7_bbfe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse := VAR_t16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;
     -- t16_MUX[uxn_opcodes_h_l961_c7_0f37] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l961_c7_0f37_cond <= VAR_t16_MUX_uxn_opcodes_h_l961_c7_0f37_cond;
     t16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue;
     t16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output := t16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l964_c7_0bed] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l964_c7_0bed] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_cond;
     result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_return_output := result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l964_c7_0bed] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_cond;
     tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue;
     tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output := tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;

     -- n16_MUX[uxn_opcodes_h_l964_c7_0bed] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l964_c7_0bed_cond <= VAR_n16_MUX_uxn_opcodes_h_l964_c7_0bed_cond;
     n16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue;
     n16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output := n16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l969_c7_8db1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l961_c7_0f37] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l969_c7_8db1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l969_c7_8db1] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l964_c7_0bed] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse := VAR_n16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l969_c7_8db1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse := VAR_t16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l961_c7_0f37] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_cond;
     tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue;
     tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output := tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;

     -- t16_MUX[uxn_opcodes_h_l953_c2_af81] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l953_c2_af81_cond <= VAR_t16_MUX_uxn_opcodes_h_l953_c2_af81_cond;
     t16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue;
     t16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l953_c2_af81_return_output := t16_MUX_uxn_opcodes_h_l953_c2_af81_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l953_c2_af81] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l964_c7_0bed] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l964_c7_0bed] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l961_c7_0f37] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l961_c7_0f37] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_cond;
     result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_return_output := result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;

     -- n16_MUX[uxn_opcodes_h_l961_c7_0f37] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l961_c7_0f37_cond <= VAR_n16_MUX_uxn_opcodes_h_l961_c7_0f37_cond;
     n16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue;
     n16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output := n16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l961_c7_0f37] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l964_c7_0bed] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse := VAR_n16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_0bed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l953_c2_af81_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l953_c2_af81] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l953_c2_af81_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l953_c2_af81_cond;
     tmp16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue;
     tmp16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l953_c2_af81_return_output := tmp16_MUX_uxn_opcodes_h_l953_c2_af81_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l953_c2_af81] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output;

     -- n16_MUX[uxn_opcodes_h_l953_c2_af81] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l953_c2_af81_cond <= VAR_n16_MUX_uxn_opcodes_h_l953_c2_af81_cond;
     n16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l953_c2_af81_iftrue;
     n16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l953_c2_af81_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l953_c2_af81_return_output := n16_MUX_uxn_opcodes_h_l953_c2_af81_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l961_c7_0f37] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l961_c7_0f37] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l961_c7_0f37] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l953_c2_af81] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_cond;
     result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_return_output := result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l953_c2_af81] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l953_c2_af81_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_0f37_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l953_c2_af81_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l953_c2_af81] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l953_c2_af81] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l953_c2_af81] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l983_l949_DUPLICATE_718c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l983_l949_DUPLICATE_718c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c2_af81_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c2_af81_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l983_l949_DUPLICATE_718c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l983_l949_DUPLICATE_718c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
