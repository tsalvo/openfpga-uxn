-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 17
entity VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_0CLK_83e31706 is
port(
 elem_val : in unsigned(7 downto 0);
 ref_toks_0 : in uint8_t_8;
 var_dim_0 : in unsigned(2 downto 0);
 return_output : out uint8_t_array_8_t);
end VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_0CLK_83e31706;
architecture arch of VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_0CLK_83e31706 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_return_output : unsigned(0 downto 0);

-- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5]
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_cond : unsigned(0 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_iftrue : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_iffalse : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_return_output : unsigned(0 downto 0);

-- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416]
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_cond : unsigned(0 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_iftrue : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_iffalse : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_return_output : unsigned(0 downto 0);

-- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c]
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_cond : unsigned(0 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_iftrue : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_iffalse : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_return_output : unsigned(0 downto 0);

-- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900]
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_cond : unsigned(0 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_iftrue : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_iffalse : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_return_output : unsigned(0 downto 0);

-- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9]
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_cond : unsigned(0 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_iftrue : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_iffalse : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_return_output : unsigned(0 downto 0);

-- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad]
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_cond : unsigned(0 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_iftrue : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_iffalse : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_return_output : unsigned(0 downto 0);

-- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de]
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_cond : unsigned(0 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_iftrue : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_iffalse : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_return_output : unsigned(0 downto 0);

-- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269]
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_cond : unsigned(0 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_iftrue : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_iffalse : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_return_output : unsigned(7 downto 0);

function CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_79ae( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return uint8_t_array_8_t is
 
  variable base : uint8_t_array_8_t; 
  variable return_output : uint8_t_array_8_t;
begin
      base.data(3) := ref_toks_0;
      base.data(2) := ref_toks_1;
      base.data(5) := ref_toks_2;
      base.data(1) := ref_toks_3;
      base.data(4) := ref_toks_4;
      base.data(7) := ref_toks_5;
      base.data(0) := ref_toks_6;
      base.data(6) := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f : entity work.BIN_OP_EQ_uint3_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_return_output);

-- rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_cond,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_iftrue,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_iffalse,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe : entity work.BIN_OP_EQ_uint3_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_return_output);

-- rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_cond,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_iftrue,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_iffalse,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163 : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_return_output);

-- rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_cond,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_iftrue,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_iffalse,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1 : entity work.BIN_OP_EQ_uint3_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_return_output);

-- rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_cond,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_iftrue,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_iffalse,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4 : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_return_output);

-- rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_cond,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_iftrue,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_iffalse,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1 : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_return_output);

-- rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_cond,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_iftrue,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_iffalse,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383 : entity work.BIN_OP_EQ_uint3_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_return_output);

-- rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_cond,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_iftrue,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_iffalse,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_return_output);

-- rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_cond,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_iftrue,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_iffalse,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 elem_val,
 ref_toks_0,
 var_dim_0,
 -- All submodule outputs
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_return_output,
 rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_return_output,
 rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_return_output,
 rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_return_output,
 rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_return_output,
 rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_return_output,
 rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_return_output,
 rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_return_output,
 rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_elem_val : unsigned(7 downto 0);
 variable VAR_ref_toks_0 : uint8_t_8;
 variable VAR_var_dim_0 : unsigned(2 downto 0);
 variable VAR_return_output : uint8_t_array_8_t;
 variable VAR_base : uint8_t_8;
 variable VAR_rv : uint8_t_array_8_t;
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_b1b1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_f5e7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_46ae_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_3895_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_7ca2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_4600_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_dac9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_cf29_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_79ae_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_2e6a_return_output : uint8_t_array_8_t;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_right := to_unsigned(7, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_elem_val := elem_val;
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_iftrue := VAR_elem_val;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_iftrue := VAR_elem_val;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_iftrue := VAR_elem_val;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_iftrue := VAR_elem_val;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_iftrue := VAR_elem_val;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_iftrue := VAR_elem_val;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_iftrue := VAR_elem_val;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_iftrue := VAR_elem_val;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_left := VAR_var_dim_0;
     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_1_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_3895] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_3895_return_output := VAR_ref_toks_0(1);

     -- CONST_REF_RD_uint8_t_uint8_t_8_5_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_46ae] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_46ae_return_output := VAR_ref_toks_0(5);

     -- CONST_REF_RD_uint8_t_uint8_t_8_3_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_b1b1] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_b1b1_return_output := VAR_ref_toks_0(3);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_6_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_cf29] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_cf29_return_output := VAR_ref_toks_0(6);

     -- CONST_REF_RD_uint8_t_uint8_t_8_7_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_4600] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_4600_return_output := VAR_ref_toks_0(7);

     -- CONST_REF_RD_uint8_t_uint8_t_8_2_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_f5e7] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_f5e7_return_output := VAR_ref_toks_0(2);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_4_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_7ca2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_7ca2_return_output := VAR_ref_toks_0(4);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_0_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_dac9] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_dac9_return_output := VAR_ref_toks_0(0);

     -- Submodule level 1
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_6a2f_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_72fe_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_f163_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_f8c1_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_8ce4_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_b7a1_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a383_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_1cab_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_dac9_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_3895_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_f5e7_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_b1b1_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_7ca2_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_46ae_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_cf29_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_4600_return_output;
     -- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416] LATENCY=0
     -- Inputs
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_cond <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_cond;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_iftrue <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_iftrue;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_iffalse <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_iffalse;
     -- Outputs
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_return_output := rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_return_output;

     -- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de] LATENCY=0
     -- Inputs
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_cond <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_cond;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_iftrue <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_iftrue;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_iffalse <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_iffalse;
     -- Outputs
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_return_output := rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_return_output;

     -- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad] LATENCY=0
     -- Inputs
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_cond <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_cond;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_iftrue <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_iftrue;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_iffalse <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_iffalse;
     -- Outputs
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_return_output := rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_return_output;

     -- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c] LATENCY=0
     -- Inputs
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_cond <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_cond;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_iftrue <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_iftrue;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_iffalse <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_iffalse;
     -- Outputs
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_return_output := rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_return_output;

     -- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5] LATENCY=0
     -- Inputs
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_cond <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_cond;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_iftrue <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_iftrue;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_iffalse <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_iffalse;
     -- Outputs
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_return_output := rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_return_output;

     -- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269] LATENCY=0
     -- Inputs
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_cond <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_cond;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_iftrue <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_iftrue;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_iffalse <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_iffalse;
     -- Outputs
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_return_output := rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_return_output;

     -- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900] LATENCY=0
     -- Inputs
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_cond <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_cond;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_iftrue <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_iftrue;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_iffalse <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_iffalse;
     -- Outputs
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_return_output := rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_return_output;

     -- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9] LATENCY=0
     -- Inputs
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_cond <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_cond;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_iftrue <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_iftrue;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_iffalse <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_iffalse;
     -- Outputs
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_return_output := rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_return_output;

     -- Submodule level 2
     -- CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_79ae[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_2e6a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_79ae_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_2e6a_return_output := CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_79ae(
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_61d5_return_output,
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3416_return_output,
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_e83c_return_output,
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_1900_return_output,
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_acd9_return_output,
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_66ad_return_output,
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_13de_return_output,
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_8269_return_output);

     -- Submodule level 3
     VAR_return_output := VAR_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_79ae_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_2e6a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
