-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity ovr_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ovr_0CLK_6d7675a8;
architecture arch of ovr_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l288_c6_24d0]
signal BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l288_c1_b3fc]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l288_c2_b0af]
signal n8_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l288_c2_b0af]
signal t8_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l288_c2_b0af]
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l288_c2_b0af]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l288_c2_b0af]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l288_c2_b0af]
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l288_c2_b0af]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l288_c2_b0af]
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l289_c3_7b34[uxn_opcodes_h_l289_c3_7b34]
signal printf_uxn_opcodes_h_l289_c3_7b34_uxn_opcodes_h_l289_c3_7b34_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l293_c11_7d54]
signal BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l293_c7_b110]
signal n8_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l293_c7_b110]
signal t8_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l293_c7_b110]
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l293_c7_b110]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l293_c7_b110]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l293_c7_b110]
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l293_c7_b110]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l293_c7_b110]
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l296_c11_d836]
signal BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l296_c7_167d]
signal n8_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l296_c7_167d]
signal t8_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l296_c7_167d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l296_c7_167d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l296_c7_167d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l296_c7_167d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l296_c7_167d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l296_c7_167d]
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l299_c11_2e35]
signal BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l299_c7_34df]
signal n8_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l299_c7_34df_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l299_c7_34df]
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l299_c7_34df]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l299_c7_34df]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l299_c7_34df]
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l299_c7_34df]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l299_c7_34df]
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l302_c30_0b84]
signal sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l307_c11_0c25]
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l307_c7_41ad]
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l307_c7_41ad]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l307_c7_41ad]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l307_c7_41ad]
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l307_c7_41ad]
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l312_c11_d871]
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l312_c7_bc76]
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l312_c7_bc76]
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l312_c7_bc76]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l312_c7_bc76]
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l316_c11_44d5]
signal BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l316_c7_4e4e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l316_c7_4e4e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5b93( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0
BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_left,
BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_right,
BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_return_output);

-- n8_MUX_uxn_opcodes_h_l288_c2_b0af
n8_MUX_uxn_opcodes_h_l288_c2_b0af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l288_c2_b0af_cond,
n8_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue,
n8_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse,
n8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output);

-- t8_MUX_uxn_opcodes_h_l288_c2_b0af
t8_MUX_uxn_opcodes_h_l288_c2_b0af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l288_c2_b0af_cond,
t8_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue,
t8_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse,
t8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af
result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_cond,
result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_return_output);

-- printf_uxn_opcodes_h_l289_c3_7b34_uxn_opcodes_h_l289_c3_7b34
printf_uxn_opcodes_h_l289_c3_7b34_uxn_opcodes_h_l289_c3_7b34 : entity work.printf_uxn_opcodes_h_l289_c3_7b34_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l289_c3_7b34_uxn_opcodes_h_l289_c3_7b34_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54
BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_left,
BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_right,
BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output);

-- n8_MUX_uxn_opcodes_h_l293_c7_b110
n8_MUX_uxn_opcodes_h_l293_c7_b110 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l293_c7_b110_cond,
n8_MUX_uxn_opcodes_h_l293_c7_b110_iftrue,
n8_MUX_uxn_opcodes_h_l293_c7_b110_iffalse,
n8_MUX_uxn_opcodes_h_l293_c7_b110_return_output);

-- t8_MUX_uxn_opcodes_h_l293_c7_b110
t8_MUX_uxn_opcodes_h_l293_c7_b110 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l293_c7_b110_cond,
t8_MUX_uxn_opcodes_h_l293_c7_b110_iftrue,
t8_MUX_uxn_opcodes_h_l293_c7_b110_iffalse,
t8_MUX_uxn_opcodes_h_l293_c7_b110_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110
result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_cond,
result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836
BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_left,
BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_right,
BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output);

-- n8_MUX_uxn_opcodes_h_l296_c7_167d
n8_MUX_uxn_opcodes_h_l296_c7_167d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l296_c7_167d_cond,
n8_MUX_uxn_opcodes_h_l296_c7_167d_iftrue,
n8_MUX_uxn_opcodes_h_l296_c7_167d_iffalse,
n8_MUX_uxn_opcodes_h_l296_c7_167d_return_output);

-- t8_MUX_uxn_opcodes_h_l296_c7_167d
t8_MUX_uxn_opcodes_h_l296_c7_167d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l296_c7_167d_cond,
t8_MUX_uxn_opcodes_h_l296_c7_167d_iftrue,
t8_MUX_uxn_opcodes_h_l296_c7_167d_iffalse,
t8_MUX_uxn_opcodes_h_l296_c7_167d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d
result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_cond,
result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35
BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_left,
BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_right,
BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_return_output);

-- n8_MUX_uxn_opcodes_h_l299_c7_34df
n8_MUX_uxn_opcodes_h_l299_c7_34df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l299_c7_34df_cond,
n8_MUX_uxn_opcodes_h_l299_c7_34df_iftrue,
n8_MUX_uxn_opcodes_h_l299_c7_34df_iffalse,
n8_MUX_uxn_opcodes_h_l299_c7_34df_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df
result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_cond,
result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_return_output);

-- sp_relative_shift_uxn_opcodes_h_l302_c30_0b84
sp_relative_shift_uxn_opcodes_h_l302_c30_0b84 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_ins,
sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_x,
sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_y,
sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25
BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_left,
BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_right,
BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad
result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_cond,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871
BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_left,
BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_right,
BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76
result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_cond,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5
BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_left,
BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_right,
BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_return_output,
 n8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output,
 t8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output,
 n8_MUX_uxn_opcodes_h_l293_c7_b110_return_output,
 t8_MUX_uxn_opcodes_h_l293_c7_b110_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output,
 n8_MUX_uxn_opcodes_h_l296_c7_167d_return_output,
 t8_MUX_uxn_opcodes_h_l296_c7_167d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_return_output,
 n8_MUX_uxn_opcodes_h_l299_c7_34df_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_return_output,
 sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l290_c3_70e4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l289_c3_7b34_uxn_opcodes_h_l289_c3_7b34_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l294_c3_a9e5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_34df_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l304_c3_2cec : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_314c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l313_c3_7e5a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_77af_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_95ec_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_2e4a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_a220_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_0191_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l296_l312_DUPLICATE_4816_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l321_l284_DUPLICATE_afb4_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_314c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_314c;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l304_c3_2cec := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l304_c3_2cec;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l313_c3_7e5a := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l313_c3_7e5a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_right := to_unsigned(6, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l294_c3_a9e5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l294_c3_a9e5;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l290_c3_70e4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l290_c3_70e4;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_b110_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_167d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_34df_iffalse := n8;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_34df_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_167d_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_b110_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_167d_iffalse := t8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l296_l312_DUPLICATE_4816 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l296_l312_DUPLICATE_4816_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_95ec LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_95ec_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_0191 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_0191_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l307_c11_0c25] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_left;
     BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_return_output := BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l316_c11_44d5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_left;
     BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_return_output := BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l293_c11_7d54] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_left;
     BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output := BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_77af LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_77af_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l302_c30_0b84] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_ins;
     sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_x <= VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_x;
     sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_y <= VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_return_output := sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_a220 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_a220_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l299_c11_2e35] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_left;
     BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_return_output := BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l312_c11_d871] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_left;
     BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_return_output := BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_2e4a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_2e4a_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l288_c6_24d0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_left;
     BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output := BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l296_c11_d836] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_left;
     BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output := BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_b0af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_b0af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_24d0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_b110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_b110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_7d54_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_167d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_167d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_d836_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_34df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_2e35_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_0c25_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_d871_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_44d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_2e4a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_2e4a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_2e4a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_2e4a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_0191_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_0191_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_0191_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_0191_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_0191_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_0191_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_95ec_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_95ec_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_95ec_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_95ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_77af_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_77af_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_77af_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_77af_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_77af_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_77af_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l296_l312_DUPLICATE_4816_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l296_l312_DUPLICATE_4816_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_a220_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_a220_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_a220_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_a220_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_0b84_return_output;
     -- n8_MUX[uxn_opcodes_h_l299_c7_34df] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l299_c7_34df_cond <= VAR_n8_MUX_uxn_opcodes_h_l299_c7_34df_cond;
     n8_MUX_uxn_opcodes_h_l299_c7_34df_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l299_c7_34df_iftrue;
     n8_MUX_uxn_opcodes_h_l299_c7_34df_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l299_c7_34df_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_34df_return_output := n8_MUX_uxn_opcodes_h_l299_c7_34df_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l316_c7_4e4e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l312_c7_bc76] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_cond;
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_return_output := result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l307_c7_41ad] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l299_c7_34df] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l312_c7_bc76] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l316_c7_4e4e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output;

     -- t8_MUX[uxn_opcodes_h_l296_c7_167d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l296_c7_167d_cond <= VAR_t8_MUX_uxn_opcodes_h_l296_c7_167d_cond;
     t8_MUX_uxn_opcodes_h_l296_c7_167d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l296_c7_167d_iftrue;
     t8_MUX_uxn_opcodes_h_l296_c7_167d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l296_c7_167d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_167d_return_output := t8_MUX_uxn_opcodes_h_l296_c7_167d_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l288_c1_b3fc] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l289_c3_7b34_uxn_opcodes_h_l289_c3_7b34_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_b3fc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_167d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l299_c7_34df_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_41ad_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_4e4e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_bc76_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_bc76_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_b110_iffalse := VAR_t8_MUX_uxn_opcodes_h_l296_c7_167d_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l296_c7_167d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output;

     -- t8_MUX[uxn_opcodes_h_l293_c7_b110] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l293_c7_b110_cond <= VAR_t8_MUX_uxn_opcodes_h_l293_c7_b110_cond;
     t8_MUX_uxn_opcodes_h_l293_c7_b110_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l293_c7_b110_iftrue;
     t8_MUX_uxn_opcodes_h_l293_c7_b110_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l293_c7_b110_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_b110_return_output := t8_MUX_uxn_opcodes_h_l293_c7_b110_return_output;

     -- printf_uxn_opcodes_h_l289_c3_7b34[uxn_opcodes_h_l289_c3_7b34] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l289_c3_7b34_uxn_opcodes_h_l289_c3_7b34_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l289_c3_7b34_uxn_opcodes_h_l289_c3_7b34_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l299_c7_34df] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l312_c7_bc76] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_return_output;

     -- n8_MUX[uxn_opcodes_h_l296_c7_167d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l296_c7_167d_cond <= VAR_n8_MUX_uxn_opcodes_h_l296_c7_167d_cond;
     n8_MUX_uxn_opcodes_h_l296_c7_167d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l296_c7_167d_iftrue;
     n8_MUX_uxn_opcodes_h_l296_c7_167d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l296_c7_167d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_167d_return_output := n8_MUX_uxn_opcodes_h_l296_c7_167d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l307_c7_41ad] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_cond;
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_return_output := result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l307_c7_41ad] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l312_c7_bc76] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_b110_iffalse := VAR_n8_MUX_uxn_opcodes_h_l296_c7_167d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_bc76_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_34df_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_bc76_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_41ad_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_41ad_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse := VAR_t8_MUX_uxn_opcodes_h_l293_c7_b110_return_output;
     -- t8_MUX[uxn_opcodes_h_l288_c2_b0af] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l288_c2_b0af_cond <= VAR_t8_MUX_uxn_opcodes_h_l288_c2_b0af_cond;
     t8_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue;
     t8_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output := t8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output;

     -- n8_MUX[uxn_opcodes_h_l293_c7_b110] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l293_c7_b110_cond <= VAR_n8_MUX_uxn_opcodes_h_l293_c7_b110_cond;
     n8_MUX_uxn_opcodes_h_l293_c7_b110_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l293_c7_b110_iftrue;
     n8_MUX_uxn_opcodes_h_l293_c7_b110_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l293_c7_b110_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_b110_return_output := n8_MUX_uxn_opcodes_h_l293_c7_b110_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l293_c7_b110] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l299_c7_34df] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_cond;
     result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_return_output := result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l299_c7_34df] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l296_c7_167d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l307_c7_41ad] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l307_c7_41ad] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse := VAR_n8_MUX_uxn_opcodes_h_l293_c7_b110_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_41ad_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_167d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_41ad_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_34df_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_34df_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l299_c7_34df] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l296_c7_167d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_return_output;

     -- n8_MUX[uxn_opcodes_h_l288_c2_b0af] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l288_c2_b0af_cond <= VAR_n8_MUX_uxn_opcodes_h_l288_c2_b0af_cond;
     n8_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue;
     n8_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output := n8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l288_c2_b0af] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l296_c7_167d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_return_output := result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l299_c7_34df] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l293_c7_b110] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l288_c2_b0af_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_34df_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_b110_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_34df_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_167d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_167d_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l296_c7_167d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l296_c7_167d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l293_c7_b110] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l293_c7_b110] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_cond;
     result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_return_output := result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l288_c2_b0af] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_167d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_167d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_b110_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_b110_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l293_c7_b110] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l293_c7_b110] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l288_c2_b0af] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_cond;
     result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_return_output := result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l288_c2_b0af] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_b110_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_b110_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l288_c2_b0af] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l288_c2_b0af] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l321_l284_DUPLICATE_afb4 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l321_l284_DUPLICATE_afb4_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5b93(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_b0af_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_b0af_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_b0af_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_b0af_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_b0af_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l321_l284_DUPLICATE_afb4_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l321_l284_DUPLICATE_afb4_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
