-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity eor_0CLK_6be78140 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor_0CLK_6be78140;
architecture arch of eor_0CLK_6be78140 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1057_c6_c782]
signal BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1057_c2_69f8]
signal n8_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1057_c2_69f8]
signal result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1057_c2_69f8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1057_c2_69f8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1057_c2_69f8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1057_c2_69f8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1057_c2_69f8]
signal t8_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1064_c11_9ce9]
signal BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1064_c7_8b14]
signal n8_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1064_c7_8b14]
signal result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1064_c7_8b14]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1064_c7_8b14]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1064_c7_8b14]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1064_c7_8b14]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1064_c7_8b14]
signal t8_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1067_c11_3617]
signal BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1067_c7_1182]
signal n8_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1067_c7_1182]
signal result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1067_c7_1182]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1067_c7_1182]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1067_c7_1182]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1067_c7_1182]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1067_c7_1182]
signal t8_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1070_c11_6dc3]
signal BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1070_c7_c2bc]
signal n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1070_c7_c2bc]
signal result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1070_c7_c2bc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1070_c7_c2bc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1070_c7_c2bc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1070_c7_c2bc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1073_c30_0214]
signal sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_return_output : signed(3 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1076_c21_205a]
signal BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_left : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_right : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1078_c11_d7db]
signal BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1078_c7_4745]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1078_c7_4745]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1078_c7_4745]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_return_output : signed(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782
BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_left,
BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_right,
BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_return_output);

-- n8_MUX_uxn_opcodes_h_l1057_c2_69f8
n8_MUX_uxn_opcodes_h_l1057_c2_69f8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1057_c2_69f8_cond,
n8_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue,
n8_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse,
n8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8
result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_cond,
result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8
result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8
result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8
result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output);

-- t8_MUX_uxn_opcodes_h_l1057_c2_69f8
t8_MUX_uxn_opcodes_h_l1057_c2_69f8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1057_c2_69f8_cond,
t8_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue,
t8_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse,
t8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9
BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_left,
BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_right,
BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_return_output);

-- n8_MUX_uxn_opcodes_h_l1064_c7_8b14
n8_MUX_uxn_opcodes_h_l1064_c7_8b14 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1064_c7_8b14_cond,
n8_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue,
n8_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse,
n8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14
result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_cond,
result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14
result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14
result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14
result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output);

-- t8_MUX_uxn_opcodes_h_l1064_c7_8b14
t8_MUX_uxn_opcodes_h_l1064_c7_8b14 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1064_c7_8b14_cond,
t8_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue,
t8_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse,
t8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617
BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_left,
BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_right,
BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_return_output);

-- n8_MUX_uxn_opcodes_h_l1067_c7_1182
n8_MUX_uxn_opcodes_h_l1067_c7_1182 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1067_c7_1182_cond,
n8_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue,
n8_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse,
n8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182
result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_cond,
result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_return_output);

-- t8_MUX_uxn_opcodes_h_l1067_c7_1182
t8_MUX_uxn_opcodes_h_l1067_c7_1182 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1067_c7_1182_cond,
t8_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue,
t8_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse,
t8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3
BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_left,
BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_right,
BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_return_output);

-- n8_MUX_uxn_opcodes_h_l1070_c7_c2bc
n8_MUX_uxn_opcodes_h_l1070_c7_c2bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond,
n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue,
n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse,
n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc
result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond,
result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc
result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc
result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc
result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1073_c30_0214
sp_relative_shift_uxn_opcodes_h_l1073_c30_0214 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_ins,
sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_x,
sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_y,
sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a
BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_left,
BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_right,
BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db
BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_left,
BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_right,
BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745
result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745
result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745
result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_return_output,
 n8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output,
 t8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_return_output,
 n8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output,
 t8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_return_output,
 n8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_return_output,
 t8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_return_output,
 n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output,
 sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1061_c3_3846 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1057_c2_69f8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1065_c3_66b0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1064_c7_8b14_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1067_c7_1182_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1075_c3_6a0c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1079_c3_00b4 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1070_l1057_l1064_l1067_DUPLICATE_130e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_e7e1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_5b16_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1070_l1064_l1078_l1067_DUPLICATE_bd88_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1070_l1067_DUPLICATE_324c_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1084_l1053_DUPLICATE_20d8_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1065_c3_66b0 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1065_c3_66b0;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1075_c3_6a0c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1075_c3_6a0c;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1061_c3_3846 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1061_c3_3846;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1079_c3_00b4 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1079_c3_00b4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1078_c11_d7db] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_left;
     BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_return_output := BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_e7e1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_e7e1_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1064_c11_9ce9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1070_c11_6dc3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_5b16 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_5b16_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1070_l1067_DUPLICATE_324c LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1070_l1067_DUPLICATE_324c_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l1073_c30_0214] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_ins;
     sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_x;
     sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_return_output := sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1070_l1057_l1064_l1067_DUPLICATE_130e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1070_l1057_l1064_l1067_DUPLICATE_130e_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1067_c11_3617] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_left;
     BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_return_output := BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_return_output;

     -- BIN_OP_XOR[uxn_opcodes_h_l1076_c21_205a] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_left;
     BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_return_output := BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1057_c6_c782] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_left;
     BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_return_output := BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1070_l1064_l1078_l1067_DUPLICATE_bd88 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1070_l1064_l1078_l1067_DUPLICATE_bd88_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1057_c2_69f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1057_c2_69f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c6_c782_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1064_c7_8b14_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1064_c7_8b14_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_9ce9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1067_c7_1182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1067_c7_1182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_3617_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1070_c11_6dc3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1078_c11_d7db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1076_c21_205a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_5b16_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_5b16_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_5b16_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_5b16_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1070_l1064_l1078_l1067_DUPLICATE_bd88_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1070_l1064_l1078_l1067_DUPLICATE_bd88_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1070_l1064_l1078_l1067_DUPLICATE_bd88_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1070_l1064_l1078_l1067_DUPLICATE_bd88_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_e7e1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_e7e1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_e7e1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1057_l1064_l1078_l1067_DUPLICATE_e7e1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1070_l1067_DUPLICATE_324c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1070_l1067_DUPLICATE_324c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1070_l1057_l1064_l1067_DUPLICATE_130e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1070_l1057_l1064_l1067_DUPLICATE_130e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1070_l1057_l1064_l1067_DUPLICATE_130e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1070_l1057_l1064_l1067_DUPLICATE_130e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1073_c30_0214_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1070_c7_c2bc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1078_c7_4745] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_return_output;

     -- n8_MUX[uxn_opcodes_h_l1070_c7_c2bc] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond <= VAR_n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond;
     n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue;
     n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output := n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1078_c7_4745] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_return_output;

     -- t8_MUX[uxn_opcodes_h_l1067_c7_1182] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1067_c7_1182_cond <= VAR_t8_MUX_uxn_opcodes_h_l1067_c7_1182_cond;
     t8_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue;
     t8_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output := t8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1070_c7_c2bc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output := result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1078_c7_4745] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1078_c7_4745_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1078_c7_4745_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1078_c7_4745_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;
     -- t8_MUX[uxn_opcodes_h_l1064_c7_8b14] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1064_c7_8b14_cond <= VAR_t8_MUX_uxn_opcodes_h_l1064_c7_8b14_cond;
     t8_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue;
     t8_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output := t8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1070_c7_c2bc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1067_c7_1182] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_return_output := result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1070_c7_c2bc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1070_c7_c2bc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1067_c7_1182] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;

     -- n8_MUX[uxn_opcodes_h_l1067_c7_1182] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1067_c7_1182_cond <= VAR_n8_MUX_uxn_opcodes_h_l1067_c7_1182_cond;
     n8_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue;
     n8_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output := n8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1070_c7_c2bc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1067_c7_1182] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1067_c7_1182] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1067_c7_1182] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;

     -- n8_MUX[uxn_opcodes_h_l1064_c7_8b14] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1064_c7_8b14_cond <= VAR_n8_MUX_uxn_opcodes_h_l1064_c7_8b14_cond;
     n8_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue;
     n8_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output := n8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1064_c7_8b14] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;

     -- t8_MUX[uxn_opcodes_h_l1057_c2_69f8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1057_c2_69f8_cond <= VAR_t8_MUX_uxn_opcodes_h_l1057_c2_69f8_cond;
     t8_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue;
     t8_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output := t8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1064_c7_8b14] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output := result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_1182_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1057_c2_69f8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output;

     -- n8_MUX[uxn_opcodes_h_l1057_c2_69f8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1057_c2_69f8_cond <= VAR_n8_MUX_uxn_opcodes_h_l1057_c2_69f8_cond;
     n8_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue;
     n8_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output := n8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1057_c2_69f8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output := result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1064_c7_8b14] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1064_c7_8b14] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1064_c7_8b14] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_8b14_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1057_c2_69f8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1057_c2_69f8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1057_c2_69f8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1084_l1053_DUPLICATE_20d8 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1084_l1053_DUPLICATE_20d8_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c2_69f8_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1084_l1053_DUPLICATE_20d8_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1084_l1053_DUPLICATE_20d8_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
