-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity sub_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub_0CLK_64d180f1;
architecture arch of sub_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2461_c6_4e55]
signal BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2461_c2_7841]
signal n8_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2461_c2_7841]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2461_c2_7841]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2461_c2_7841]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2461_c2_7841]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2461_c2_7841]
signal result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2461_c2_7841]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2461_c2_7841]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2461_c2_7841]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2461_c2_7841]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2461_c2_7841]
signal t8_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2474_c11_1edd]
signal BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2474_c7_0cff]
signal n8_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2474_c7_0cff]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2474_c7_0cff]
signal result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2474_c7_0cff]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2474_c7_0cff]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2474_c7_0cff]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2474_c7_0cff]
signal t8_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2477_c11_320c]
signal BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2477_c7_3794]
signal n8_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2477_c7_3794]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2477_c7_3794]
signal result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2477_c7_3794]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2477_c7_3794]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2477_c7_3794]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2477_c7_3794]
signal t8_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2480_c11_7326]
signal BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2480_c7_6586]
signal n8_MUX_uxn_opcodes_h_l2480_c7_6586_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2480_c7_6586_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2480_c7_6586]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2480_c7_6586]
signal result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2480_c7_6586]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2480_c7_6586]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2480_c7_6586]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2482_c30_c549]
signal sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_return_output : signed(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2485_c21_8ed9]
signal BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_opc_done := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55
BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_left,
BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_right,
BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output);

-- n8_MUX_uxn_opcodes_h_l2461_c2_7841
n8_MUX_uxn_opcodes_h_l2461_c2_7841 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2461_c2_7841_cond,
n8_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue,
n8_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse,
n8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_cond,
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_return_output);

-- t8_MUX_uxn_opcodes_h_l2461_c2_7841
t8_MUX_uxn_opcodes_h_l2461_c2_7841 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2461_c2_7841_cond,
t8_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue,
t8_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse,
t8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd
BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_left,
BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_right,
BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_return_output);

-- n8_MUX_uxn_opcodes_h_l2474_c7_0cff
n8_MUX_uxn_opcodes_h_l2474_c7_0cff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2474_c7_0cff_cond,
n8_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue,
n8_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse,
n8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_cond,
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output);

-- t8_MUX_uxn_opcodes_h_l2474_c7_0cff
t8_MUX_uxn_opcodes_h_l2474_c7_0cff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2474_c7_0cff_cond,
t8_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue,
t8_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse,
t8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c
BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_left,
BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_right,
BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_return_output);

-- n8_MUX_uxn_opcodes_h_l2477_c7_3794
n8_MUX_uxn_opcodes_h_l2477_c7_3794 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2477_c7_3794_cond,
n8_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue,
n8_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse,
n8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_cond,
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_return_output);

-- t8_MUX_uxn_opcodes_h_l2477_c7_3794
t8_MUX_uxn_opcodes_h_l2477_c7_3794 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2477_c7_3794_cond,
t8_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue,
t8_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse,
t8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326
BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_left,
BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_right,
BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_return_output);

-- n8_MUX_uxn_opcodes_h_l2480_c7_6586
n8_MUX_uxn_opcodes_h_l2480_c7_6586 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2480_c7_6586_cond,
n8_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue,
n8_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse,
n8_MUX_uxn_opcodes_h_l2480_c7_6586_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_cond,
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2482_c30_c549
sp_relative_shift_uxn_opcodes_h_l2482_c30_c549 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_ins,
sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_x,
sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_y,
sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9
BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_left,
BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_right,
BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output,
 n8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
 t8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_return_output,
 n8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output,
 t8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_return_output,
 n8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_return_output,
 t8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_return_output,
 n8_MUX_uxn_opcodes_h_l2480_c7_6586_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_return_output,
 sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2466_c3_8ef6 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2471_c3_041e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2461_c2_7841_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2475_c3_1aa1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2474_c7_0cff_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2480_c7_6586_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2477_c7_3794_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2480_c7_6586_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2484_c3_7531 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_f2cc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_8d5d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_46e6_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_9b0b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2477_l2480_DUPLICATE_5e3c_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2457_l2489_DUPLICATE_b87c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2471_c3_041e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2471_c3_041e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_right := to_unsigned(2, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2475_c3_1aa1 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2475_c3_1aa1;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2466_c3_8ef6 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2466_c3_8ef6;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2484_c3_7531 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2484_c3_7531;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_8d5d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_8d5d_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_f2cc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_f2cc_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2477_c11_320c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_return_output;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2485_c21_8ed9] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2461_c2_7841_return_output := result.is_ram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2461_c2_7841_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2461_c6_4e55] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_left;
     BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output := BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2480_c11_7326] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_left;
     BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_return_output := BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_9b0b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_9b0b_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l2482_c30_c549] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_ins;
     sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_x;
     sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_return_output := sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2474_c11_1edd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2461_c2_7841_return_output := result.is_vram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2461_c2_7841_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2477_l2480_DUPLICATE_5e3c LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2477_l2480_DUPLICATE_5e3c_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_46e6 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_46e6_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2461_c2_7841_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2461_c2_7841_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_4e55_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2474_c7_0cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2474_c7_0cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_1edd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2477_c7_3794_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2477_c7_3794_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_320c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2480_c7_6586_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_7326_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_8ed9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_46e6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_46e6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_46e6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_9b0b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_9b0b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_9b0b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_8d5d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_8d5d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2477_l2480_l2474_DUPLICATE_8d5d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2477_l2480_DUPLICATE_5e3c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2477_l2480_DUPLICATE_5e3c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_f2cc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_f2cc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_f2cc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2477_l2461_l2480_l2474_DUPLICATE_f2cc_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2461_c2_7841_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2461_c2_7841_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2461_c2_7841_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2461_c2_7841_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_c549_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2480_c7_6586] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2480_c7_6586] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_return_output;

     -- n8_MUX[uxn_opcodes_h_l2480_c7_6586] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2480_c7_6586_cond <= VAR_n8_MUX_uxn_opcodes_h_l2480_c7_6586_cond;
     n8_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue;
     n8_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2480_c7_6586_return_output := n8_MUX_uxn_opcodes_h_l2480_c7_6586_return_output;

     -- t8_MUX[uxn_opcodes_h_l2477_c7_3794] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2477_c7_3794_cond <= VAR_t8_MUX_uxn_opcodes_h_l2477_c7_3794_cond;
     t8_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue;
     t8_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output := t8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2480_c7_6586] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2480_c7_6586] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_return_output := result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2480_c7_6586] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2480_c7_6586_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_6586_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_6586_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_6586_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_6586_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_6586_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;
     -- t8_MUX[uxn_opcodes_h_l2474_c7_0cff] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2474_c7_0cff_cond <= VAR_t8_MUX_uxn_opcodes_h_l2474_c7_0cff_cond;
     t8_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue;
     t8_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output := t8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2477_c7_3794] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_return_output := result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2477_c7_3794] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2477_c7_3794] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2477_c7_3794] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;

     -- n8_MUX[uxn_opcodes_h_l2477_c7_3794] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2477_c7_3794_cond <= VAR_n8_MUX_uxn_opcodes_h_l2477_c7_3794_cond;
     n8_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue;
     n8_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output := n8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2477_c7_3794] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_3794_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2474_c7_0cff] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2474_c7_0cff] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2474_c7_0cff] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;

     -- n8_MUX[uxn_opcodes_h_l2474_c7_0cff] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2474_c7_0cff_cond <= VAR_n8_MUX_uxn_opcodes_h_l2474_c7_0cff_cond;
     n8_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue;
     n8_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output := n8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2474_c7_0cff] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;

     -- t8_MUX[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2461_c2_7841_cond <= VAR_t8_MUX_uxn_opcodes_h_l2461_c2_7841_cond;
     t8_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue;
     t8_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output := t8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2474_c7_0cff] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output := result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_0cff_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output;

     -- n8_MUX[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2461_c2_7841_cond <= VAR_n8_MUX_uxn_opcodes_h_l2461_c2_7841_cond;
     n8_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue;
     n8_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output := n8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_return_output := result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2461_c2_7841] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2461_c2_7841_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2457_l2489_DUPLICATE_b87c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2457_l2489_DUPLICATE_b87c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_7841_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_7841_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2457_l2489_DUPLICATE_b87c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2457_l2489_DUPLICATE_b87c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
