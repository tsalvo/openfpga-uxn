-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 30
entity lit_0CLK_ac9ce6a4 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lit_0CLK_ac9ce6a4;
architecture arch of lit_0CLK_ac9ce6a4 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l181_c6_612b]
signal BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l181_c1_1835]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l181_c2_94c9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l181_c2_94c9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l181_c2_94c9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l181_c2_94c9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l181_c2_94c9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l181_c2_94c9]
signal result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l181_c2_94c9]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l181_c2_94c9]
signal result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l182_c3_2525[uxn_opcodes_h_l182_c3_2525]
signal printf_uxn_opcodes_h_l182_c3_2525_uxn_opcodes_h_l182_c3_2525_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l188_c11_5ce5]
signal BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l188_c7_6c4d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l188_c7_6c4d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l188_c7_6c4d]
signal result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l188_c7_6c4d]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l188_c7_6c4d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l188_c7_6c4d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l188_c7_6c4d]
signal result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l191_c22_7f09]
signal BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l193_c11_6c03]
signal BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l193_c7_a920]
signal result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l193_c7_a920]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l193_c7_a920]
signal result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l193_c7_a920]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l193_c7_a920]
signal result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l199_c11_14d0]
signal BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l199_c7_c63d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l199_c7_c63d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_219b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : signed;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.sp_relative_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.u8_value := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.u16_value := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b
BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_left,
BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_right,
BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9
result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9
result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9
result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9
result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9
result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_cond,
result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9
result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9
result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_cond,
result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output);

-- printf_uxn_opcodes_h_l182_c3_2525_uxn_opcodes_h_l182_c3_2525
printf_uxn_opcodes_h_l182_c3_2525_uxn_opcodes_h_l182_c3_2525 : entity work.printf_uxn_opcodes_h_l182_c3_2525_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l182_c3_2525_uxn_opcodes_h_l182_c3_2525_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5
BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_left,
BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_right,
BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d
result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d
result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_cond,
result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d
result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d
result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d
result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d
result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_cond,
result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09
BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09 : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_left,
BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_right,
BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03
BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_left,
BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_right,
BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920
result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920
result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_cond,
result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920
result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920
result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0
BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_left,
BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_right,
BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d
result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d
result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 previous_ram_read,
 -- Registers
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l184_c3_04df : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l181_c2_94c9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l182_c3_2525_uxn_opcodes_h_l182_c3_2525_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l191_c3_5d5b : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l188_c7_6c4d_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l196_c3_6f0f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l193_l181_l188_DUPLICATE_8fc2_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l181_l199_l188_DUPLICATE_8625_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l193_l181_l188_DUPLICATE_013e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l193_l181_DUPLICATE_d78e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l193_l199_l188_DUPLICATE_b20e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_219b_uxn_opcodes_h_l177_l204_DUPLICATE_644e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_sp_relative_shift_uxn_opcodes_h_l184_c3_04df := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l184_c3_04df;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l196_c3_6f0f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l196_c3_6f0f;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_left := VAR_pc;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_iftrue := VAR_previous_ram_read;
     -- BIN_OP_EQ[uxn_opcodes_h_l188_c11_5ce5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_left;
     BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_return_output := BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l193_c11_6c03] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_left;
     BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_return_output := BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_return_output;

     -- result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d[uxn_opcodes_h_l188_c7_6c4d] LATENCY=0
     VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l188_c7_6c4d_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l181_c6_612b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_left;
     BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output := BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l193_l199_l188_DUPLICATE_b20e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l193_l199_l188_DUPLICATE_b20e_return_output := result.is_opc_done;

     -- BIN_OP_PLUS[uxn_opcodes_h_l191_c22_7f09] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_left;
     BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_return_output := BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l193_l181_DUPLICATE_d78e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l193_l181_DUPLICATE_d78e_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l193_l181_l188_DUPLICATE_013e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l193_l181_l188_DUPLICATE_013e_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l181_l199_l188_DUPLICATE_8625 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l181_l199_l188_DUPLICATE_8625_return_output := result.is_stack_write;

     -- result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d[uxn_opcodes_h_l188_c7_6c4d] LATENCY=0
     VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l188_c7_6c4d_return_output := result.is_sp_shift;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l181_c2_94c9] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l181_c2_94c9_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l199_c11_14d0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_left;
     BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_return_output := BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l193_l181_l188_DUPLICATE_8fc2 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l193_l181_l188_DUPLICATE_8fc2_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l181_c6_612b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l188_c11_5ce5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l193_c11_6c03_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l199_c11_14d0_return_output;
     VAR_result_u16_value_uxn_opcodes_h_l191_c3_5d5b := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l191_c22_7f09_return_output, 16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l193_l199_l188_DUPLICATE_b20e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l193_l199_l188_DUPLICATE_b20e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l193_l199_l188_DUPLICATE_b20e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l193_l181_DUPLICATE_d78e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l193_l181_DUPLICATE_d78e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l181_l199_l188_DUPLICATE_8625_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l181_l199_l188_DUPLICATE_8625_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l181_l199_l188_DUPLICATE_8625_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l193_l181_l188_DUPLICATE_8fc2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l193_l181_l188_DUPLICATE_8fc2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l193_l181_l188_DUPLICATE_8fc2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l193_l181_l188_DUPLICATE_013e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l193_l181_l188_DUPLICATE_013e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l193_l181_l188_DUPLICATE_013e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse := VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l188_c7_6c4d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l181_c2_94c9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse := VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l188_c7_6c4d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue := VAR_result_u16_value_uxn_opcodes_h_l191_c3_5d5b;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l181_c1_1835] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l188_c7_6c4d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l181_c2_94c9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l188_c7_6c4d] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_cond;
     result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output := result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l193_c7_a920] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_cond;
     result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_return_output := result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l193_c7_a920] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l199_c7_c63d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l199_c7_c63d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l193_c7_a920] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l182_c3_2525_uxn_opcodes_h_l182_c3_2525_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l181_c1_1835_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l199_c7_c63d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l193_c7_a920_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l199_c7_c63d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l193_c7_a920_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l193_c7_a920_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l188_c7_6c4d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output := result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l181_c2_94c9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output := result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l181_c2_94c9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l193_c7_a920] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_return_output;

     -- printf_uxn_opcodes_h_l182_c3_2525[uxn_opcodes_h_l182_c3_2525] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l182_c3_2525_uxn_opcodes_h_l182_c3_2525_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l182_c3_2525_uxn_opcodes_h_l182_c3_2525_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l188_c7_6c4d] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l193_c7_a920] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l188_c7_6c4d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l193_c7_a920_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l193_c7_a920_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l181_c2_94c9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output := result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l188_c7_6c4d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l188_c7_6c4d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l181_c2_94c9] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l181_c2_94c9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l188_c7_6c4d_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l181_c2_94c9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l181_c2_94c9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_return_output;

     -- Submodule level 5
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_219b_uxn_opcodes_h_l177_l204_DUPLICATE_644e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_219b_uxn_opcodes_h_l177_l204_DUPLICATE_644e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_219b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l181_c2_94c9_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l181_c2_94c9_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_219b_uxn_opcodes_h_l177_l204_DUPLICATE_644e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_219b_uxn_opcodes_h_l177_l204_DUPLICATE_644e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
