-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity sta_0CLK_bce25fe8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sta_0CLK_bce25fe8;
architecture arch of sta_0CLK_bce25fe8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2315_c6_f05f]
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2315_c2_4438]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2315_c2_4438]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2315_c2_4438]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2315_c2_4438]
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2315_c2_4438]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2315_c2_4438]
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2315_c2_4438]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2315_c2_4438]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2315_c2_4438]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2315_c2_4438]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2315_c2_4438]
signal n8_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2315_c2_4438]
signal t16_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2328_c11_5f5e]
signal BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2328_c7_a767]
signal result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2328_c7_a767]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2328_c7_a767]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2328_c7_a767]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2328_c7_a767]
signal result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2328_c7_a767]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2328_c7_a767]
signal n8_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2328_c7_a767]
signal t16_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2331_c11_6462]
signal BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2331_c7_5d91]
signal result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2331_c7_5d91]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2331_c7_5d91]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2331_c7_5d91]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2331_c7_5d91]
signal result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2331_c7_5d91]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2331_c7_5d91]
signal n8_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2331_c7_5d91]
signal t16_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2333_c3_96b3]
signal CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2336_c11_c7c0]
signal BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2336_c7_e0ea]
signal result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2336_c7_e0ea]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2336_c7_e0ea]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2336_c7_e0ea]
signal result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2336_c7_e0ea]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2336_c7_e0ea]
signal n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2336_c7_e0ea]
signal t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2337_c3_7709]
signal BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2339_c11_df3a]
signal BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2339_c7_3767]
signal result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2339_c7_3767]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2339_c7_3767]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2339_c7_3767]
signal result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2339_c7_3767]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2339_c7_3767]
signal n8_MUX_uxn_opcodes_h_l2339_c7_3767_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2339_c7_3767_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2341_c30_f96a]
signal sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_return_output : signed(3 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_775a( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.u16_value := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;
      base.is_ram_write := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f
BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_left,
BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_right,
BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438
result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438
result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_cond,
result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438
result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_cond,
result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438
result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output);

-- n8_MUX_uxn_opcodes_h_l2315_c2_4438
n8_MUX_uxn_opcodes_h_l2315_c2_4438 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2315_c2_4438_cond,
n8_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue,
n8_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse,
n8_MUX_uxn_opcodes_h_l2315_c2_4438_return_output);

-- t16_MUX_uxn_opcodes_h_l2315_c2_4438
t16_MUX_uxn_opcodes_h_l2315_c2_4438 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2315_c2_4438_cond,
t16_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue,
t16_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse,
t16_MUX_uxn_opcodes_h_l2315_c2_4438_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e
BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_left,
BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_right,
BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767
result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_cond,
result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767
result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767
result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767
result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_cond,
result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767
result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_return_output);

-- n8_MUX_uxn_opcodes_h_l2328_c7_a767
n8_MUX_uxn_opcodes_h_l2328_c7_a767 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2328_c7_a767_cond,
n8_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue,
n8_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse,
n8_MUX_uxn_opcodes_h_l2328_c7_a767_return_output);

-- t16_MUX_uxn_opcodes_h_l2328_c7_a767
t16_MUX_uxn_opcodes_h_l2328_c7_a767 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2328_c7_a767_cond,
t16_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue,
t16_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse,
t16_MUX_uxn_opcodes_h_l2328_c7_a767_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462
BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_left,
BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_right,
BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91
result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_cond,
result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91
result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91
result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_cond,
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output);

-- n8_MUX_uxn_opcodes_h_l2331_c7_5d91
n8_MUX_uxn_opcodes_h_l2331_c7_5d91 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2331_c7_5d91_cond,
n8_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue,
n8_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse,
n8_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output);

-- t16_MUX_uxn_opcodes_h_l2331_c7_5d91
t16_MUX_uxn_opcodes_h_l2331_c7_5d91 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2331_c7_5d91_cond,
t16_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue,
t16_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse,
t16_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3
CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3_x,
CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0
BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_left,
BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_right,
BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea
result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond,
result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea
result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea
result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond,
result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output);

-- n8_MUX_uxn_opcodes_h_l2336_c7_e0ea
n8_MUX_uxn_opcodes_h_l2336_c7_e0ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond,
n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue,
n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse,
n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output);

-- t16_MUX_uxn_opcodes_h_l2336_c7_e0ea
t16_MUX_uxn_opcodes_h_l2336_c7_e0ea : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond,
t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue,
t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse,
t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709
BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_left,
BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_right,
BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a
BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_left,
BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_right,
BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767
result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_cond,
result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767
result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_cond,
result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_return_output);

-- n8_MUX_uxn_opcodes_h_l2339_c7_3767
n8_MUX_uxn_opcodes_h_l2339_c7_3767 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2339_c7_3767_cond,
n8_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue,
n8_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse,
n8_MUX_uxn_opcodes_h_l2339_c7_3767_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a
sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_ins,
sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_x,
sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_y,
sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
 n8_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
 t16_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_return_output,
 n8_MUX_uxn_opcodes_h_l2328_c7_a767_return_output,
 t16_MUX_uxn_opcodes_h_l2328_c7_a767_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output,
 n8_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output,
 t16_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output,
 CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output,
 n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output,
 t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_return_output,
 n8_MUX_uxn_opcodes_h_l2339_c7_3767_return_output,
 sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2320_c3_058b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2325_c3_f39c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2328_c7_a767_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c2_4438_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c2_4438_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2329_c3_6973 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2328_c7_a767_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2334_c3_b48a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2331_c7_5d91_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2331_c7_5d91_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2339_c7_3767_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2339_c7_3767_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_9680_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_28c3_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_d3bc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_85dd_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0d8d_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2332_l2337_DUPLICATE_c99a_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_775a_uxn_opcodes_h_l2348_l2310_DUPLICATE_d4df_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2334_c3_b48a := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2334_c3_b48a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_right := to_unsigned(2, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_right := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_right := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2329_c3_6973 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2329_c3_6973;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2320_c3_058b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2320_c3_058b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_y := resize(to_signed(-3, 3), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2325_c3_f39c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2325_c3_f39c;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_left := t16;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse := t16;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_85dd LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_85dd_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2339_c11_df3a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2336_c11_c7c0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2341_c30_f96a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_ins;
     sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_x;
     sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_return_output := sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2315_c2_4438_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_28c3 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_28c3_return_output := result.u16_value;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2332_l2337_DUPLICATE_c99a LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2332_l2337_DUPLICATE_c99a_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2331_c7_5d91] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2331_c7_5d91_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_9680 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_9680_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2331_c11_6462] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_left;
     BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output := BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_d3bc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_d3bc_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0d8d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0d8d_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2328_c11_5f5e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2315_c2_4438_return_output := result.is_stack_index_flipped;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2315_c2_4438_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2315_c6_f05f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2315_c2_4438_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2315_c2_4438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c2_4438_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_f05f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2328_c7_a767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2328_c7_a767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_5f5e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2331_c7_5d91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2331_c7_5d91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_6462_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_c7c0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2339_c7_3767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_df3a_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2332_l2337_DUPLICATE_c99a_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2332_l2337_DUPLICATE_c99a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_85dd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_85dd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_85dd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_85dd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_28c3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_28c3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_28c3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_28c3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_28c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0d8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0d8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0d8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0d8d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_d3bc_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_d3bc_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_d3bc_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_d3bc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_9680_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_9680_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_9680_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_9680_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2339_l2336_l2331_l2328_l2315_DUPLICATE_9680_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2315_c2_4438_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2315_c2_4438_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2315_c2_4438_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2315_c2_4438_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2331_c7_5d91_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_f96a_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;

     -- n8_MUX[uxn_opcodes_h_l2339_c7_3767] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2339_c7_3767_cond <= VAR_n8_MUX_uxn_opcodes_h_l2339_c7_3767_cond;
     n8_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue;
     n8_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2339_c7_3767_return_output := n8_MUX_uxn_opcodes_h_l2339_c7_3767_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2339_c7_3767] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2331_c7_5d91] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l2333_c3_96b3] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3_return_output := CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2339_c7_3767] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output := result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2339_c7_3767] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output := result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2339_c7_3767] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2337_c3_7709] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_left;
     BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_return_output := BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2339_c7_3767] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_7709_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2333_c3_96b3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2339_c7_3767_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_3767_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_3767_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_3767_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_3767_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2336_c7_e0ea] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2336_c7_e0ea] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2336_c7_e0ea] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;

     -- n8_MUX[uxn_opcodes_h_l2336_c7_e0ea] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond <= VAR_n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond;
     n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue;
     n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output := n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2336_c7_e0ea] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output := result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2336_c7_e0ea] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output := result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;

     -- t16_MUX[uxn_opcodes_h_l2336_c7_e0ea] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond <= VAR_t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_cond;
     t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_iftrue;
     t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output := t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2328_c7_a767] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2336_c7_e0ea_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2331_c7_5d91] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output := result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2331_c7_5d91] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2331_c7_5d91] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;

     -- n8_MUX[uxn_opcodes_h_l2331_c7_5d91] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2331_c7_5d91_cond <= VAR_n8_MUX_uxn_opcodes_h_l2331_c7_5d91_cond;
     n8_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue;
     n8_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output := n8_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;

     -- t16_MUX[uxn_opcodes_h_l2331_c7_5d91] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2331_c7_5d91_cond <= VAR_t16_MUX_uxn_opcodes_h_l2331_c7_5d91_cond;
     t16_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue;
     t16_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output := t16_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2331_c7_5d91] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output := result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2331_c7_5d91] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2331_c7_5d91_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l2328_c7_a767] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;

     -- n8_MUX[uxn_opcodes_h_l2328_c7_a767] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2328_c7_a767_cond <= VAR_n8_MUX_uxn_opcodes_h_l2328_c7_a767_cond;
     n8_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue;
     n8_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2328_c7_a767_return_output := n8_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2328_c7_a767] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2328_c7_a767] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output := result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;

     -- t16_MUX[uxn_opcodes_h_l2328_c7_a767] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2328_c7_a767_cond <= VAR_t16_MUX_uxn_opcodes_h_l2328_c7_a767_cond;
     t16_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue;
     t16_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2328_c7_a767_return_output := t16_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2328_c7_a767] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2328_c7_a767] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output := result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2328_c7_a767_return_output;
     -- t16_MUX[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2315_c2_4438_cond <= VAR_t16_MUX_uxn_opcodes_h_l2315_c2_4438_cond;
     t16_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue;
     t16_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2315_c2_4438_return_output := t16_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output := result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;

     -- n8_MUX[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2315_c2_4438_cond <= VAR_n8_MUX_uxn_opcodes_h_l2315_c2_4438_cond;
     n8_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue;
     n8_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2315_c2_4438_return_output := n8_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2315_c2_4438] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output := result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2315_c2_4438_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_775a_uxn_opcodes_h_l2348_l2310_DUPLICATE_d4df LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_775a_uxn_opcodes_h_l2348_l2310_DUPLICATE_d4df_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_775a(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_4438_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_4438_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_775a_uxn_opcodes_h_l2348_l2310_DUPLICATE_d4df_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_775a_uxn_opcodes_h_l2348_l2310_DUPLICATE_d4df_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
