-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity ldz_0CLK_b128164d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_b128164d;
architecture arch of ldz_0CLK_b128164d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1460_c6_5bc8]
signal BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1460_c2_bc2c]
signal t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1460_c2_bc2c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1460_c2_bc2c]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1460_c2_bc2c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1460_c2_bc2c]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1460_c2_bc2c]
signal result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1460_c2_bc2c]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1460_c2_bc2c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1460_c2_bc2c]
signal result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1460_c2_bc2c]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1460_c2_bc2c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1460_c2_bc2c]
signal tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1473_c11_607d]
signal BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1473_c7_30e8]
signal t8_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1473_c7_30e8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1473_c7_30e8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1473_c7_30e8]
signal result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1473_c7_30e8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1473_c7_30e8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1473_c7_30e8]
signal result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1473_c7_30e8]
signal tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1476_c11_a2c1]
signal BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1476_c7_e1da]
signal t8_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1476_c7_e1da]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1476_c7_e1da]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1476_c7_e1da]
signal result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1476_c7_e1da]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1476_c7_e1da]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1476_c7_e1da]
signal result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1476_c7_e1da]
signal tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1478_c30_9aff]
signal sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1481_c11_25da]
signal BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1481_c7_85a3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1481_c7_85a3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1481_c7_85a3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1481_c7_85a3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1481_c7_85a3]
signal result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1481_c7_85a3]
signal tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1484_c11_e028]
signal BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1484_c7_f155]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1484_c7_f155]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1484_c7_f155]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1484_c7_f155]
signal result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1484_c7_f155]
signal tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_return_output : unsigned(7 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.u16_value := ref_toks_8;
      base.is_pc_updated := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8
BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_left,
BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_right,
BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output);

-- t8_MUX_uxn_opcodes_h_l1460_c2_bc2c
t8_MUX_uxn_opcodes_h_l1460_c2_bc2c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond,
t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue,
t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse,
t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c
result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c
result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c
result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c
result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c
result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond,
result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c
result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c
result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c
tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond,
tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue,
tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse,
tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d
BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_left,
BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_right,
BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output);

-- t8_MUX_uxn_opcodes_h_l1473_c7_30e8
t8_MUX_uxn_opcodes_h_l1473_c7_30e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1473_c7_30e8_cond,
t8_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue,
t8_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse,
t8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8
result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8
result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_cond,
result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8
result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8
result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8
result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_cond,
result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8
tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_cond,
tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue,
tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse,
tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1
BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_left,
BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_right,
BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output);

-- t8_MUX_uxn_opcodes_h_l1476_c7_e1da
t8_MUX_uxn_opcodes_h_l1476_c7_e1da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1476_c7_e1da_cond,
t8_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue,
t8_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse,
t8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da
result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da
result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_cond,
result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da
result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da
result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da
result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_cond,
result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da
tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_cond,
tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue,
tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse,
tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff
sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_ins,
sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_x,
sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_y,
sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da
BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_left,
BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_right,
BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3
result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3
result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3
result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3
result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_cond,
result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3
tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_cond,
tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue,
tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse,
tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028
BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_left,
BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_right,
BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155
result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155
result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155
result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_cond,
result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1484_c7_f155
tmp8_MUX_uxn_opcodes_h_l1484_c7_f155 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_cond,
tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue,
tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse,
tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output,
 t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
 tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output,
 t8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output,
 tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output,
 t8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output,
 tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output,
 sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output,
 tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_return_output,
 tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1465_c3_6a00 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1470_c3_f31a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1474_c3_06ba : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1479_c22_3b67_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1482_c3_5d1b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1487_c3_0991 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1484_l1481_l1476_l1473_l1460_DUPLICATE_1862_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1473_l1476_l1460_DUPLICATE_9f44_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_0816_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1473_l1481_DUPLICATE_874c_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_a767_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1484_l1476_l1481_DUPLICATE_3b9d_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1456_l1492_DUPLICATE_0d5a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_right := to_unsigned(2, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1487_c3_0991 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1487_c3_0991;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1465_c3_6a00 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1465_c3_6a00;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_right := to_unsigned(3, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1482_c3_5d1b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1482_c3_5d1b;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1470_c3_f31a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1470_c3_f31a;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1474_c3_06ba := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1474_c3_06ba;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse := tmp8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_a767 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_a767_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_0816 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_0816_return_output := result.is_stack_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1460_c2_bc2c_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l1478_c30_9aff] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_ins;
     sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_x;
     sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_return_output := sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1460_c2_bc2c_return_output := result.is_vram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1460_c2_bc2c_return_output := result.is_pc_updated;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1460_c2_bc2c_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1460_c6_5bc8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1473_l1476_l1460_DUPLICATE_9f44 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1473_l1476_l1460_DUPLICATE_9f44_return_output := result.u16_value;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1479_c22_3b67] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1479_c22_3b67_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1473_l1481_DUPLICATE_874c LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1473_l1481_DUPLICATE_874c_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1484_l1476_l1481_DUPLICATE_3b9d LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1484_l1476_l1481_DUPLICATE_3b9d_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1484_c11_e028] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_left;
     BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_return_output := BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1481_c11_25da] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_left;
     BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_return_output := BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1473_c11_607d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1484_l1481_l1476_l1473_l1460_DUPLICATE_1862 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1484_l1481_l1476_l1473_l1460_DUPLICATE_1862_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1476_c11_a2c1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c6_5bc8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1473_c7_30e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1473_c11_607d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1476_c7_e1da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c11_a2c1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1481_c11_25da_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1484_c11_e028_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1479_c22_3b67_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1473_l1481_DUPLICATE_874c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1473_l1481_DUPLICATE_874c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1473_l1476_l1460_DUPLICATE_9f44_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1473_l1476_l1460_DUPLICATE_9f44_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1473_l1476_l1460_DUPLICATE_9f44_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_a767_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_a767_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_a767_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_a767_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_0816_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_0816_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_0816_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1473_l1484_l1476_l1481_DUPLICATE_0816_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1484_l1476_l1481_DUPLICATE_3b9d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1484_l1476_l1481_DUPLICATE_3b9d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1484_l1476_l1481_DUPLICATE_3b9d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1484_l1481_l1476_l1473_l1460_DUPLICATE_1862_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1484_l1481_l1476_l1473_l1460_DUPLICATE_1862_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1484_l1481_l1476_l1473_l1460_DUPLICATE_1862_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1484_l1481_l1476_l1473_l1460_DUPLICATE_1862_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1484_l1481_l1476_l1473_l1460_DUPLICATE_1862_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1460_c2_bc2c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1460_c2_bc2c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1460_c2_bc2c_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1460_c2_bc2c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1478_c30_9aff_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1484_c7_f155] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_return_output := result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_return_output;

     -- t8_MUX[uxn_opcodes_h_l1476_c7_e1da] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1476_c7_e1da_cond <= VAR_t8_MUX_uxn_opcodes_h_l1476_c7_e1da_cond;
     t8_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue;
     t8_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output := t8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1476_c7_e1da] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output := result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1481_c7_85a3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1484_c7_f155] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1484_c7_f155] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_cond;
     tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_return_output := tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1484_c7_f155] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1484_c7_f155] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1484_c7_f155_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1484_c7_f155_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1484_c7_f155_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1484_c7_f155_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1484_c7_f155_return_output;
     -- t8_MUX[uxn_opcodes_h_l1473_c7_30e8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1473_c7_30e8_cond <= VAR_t8_MUX_uxn_opcodes_h_l1473_c7_30e8_cond;
     t8_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue;
     t8_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output := t8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1481_c7_85a3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1481_c7_85a3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1481_c7_85a3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1481_c7_85a3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output := result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1476_c7_e1da] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1481_c7_85a3] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_cond;
     tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output := tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1473_c7_30e8] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output := result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1481_c7_85a3_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1476_c7_e1da] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1476_c7_e1da] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output := result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1476_c7_e1da] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1476_c7_e1da] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1473_c7_30e8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;

     -- t8_MUX[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond <= VAR_t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond;
     t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue;
     t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output := t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output := result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1476_c7_e1da] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_cond;
     tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output := tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1476_c7_e1da_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1473_c7_30e8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1473_c7_30e8] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_cond;
     tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output := tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1473_c7_30e8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1473_c7_30e8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1473_c7_30e8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output := result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1473_c7_30e8_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond;
     tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output := tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1460_c2_bc2c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;

     -- Submodule level 6
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1456_l1492_DUPLICATE_0d5a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1456_l1492_DUPLICATE_0d5a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c2_bc2c_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1456_l1492_DUPLICATE_0d5a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1456_l1492_DUPLICATE_0d5a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
