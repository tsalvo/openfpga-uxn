-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 43
entity inc_0CLK_66ba3dc0 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc_0CLK_66ba3dc0;
architecture arch of inc_0CLK_66ba3dc0 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1332_c6_b074]
signal BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1332_c1_5c08]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1332_c2_0ed7]
signal t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1332_c2_0ed7]
signal result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1332_c2_0ed7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1332_c2_0ed7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1332_c2_0ed7]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1332_c2_0ed7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1332_c2_0ed7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1332_c2_0ed7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l1333_c3_da23[uxn_opcodes_h_l1333_c3_da23]
signal printf_uxn_opcodes_h_l1333_c3_da23_uxn_opcodes_h_l1333_c3_da23_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1338_c11_3b61]
signal BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1338_c7_8e08]
signal t8_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1338_c7_8e08]
signal result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1338_c7_8e08]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1338_c7_8e08]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1338_c7_8e08]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1338_c7_8e08]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1338_c7_8e08]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1338_c7_8e08]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1341_c11_0434]
signal BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1341_c7_4d29]
signal t8_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1341_c7_4d29]
signal result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1341_c7_4d29]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1341_c7_4d29]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1341_c7_4d29]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1341_c7_4d29]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1341_c7_4d29]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1341_c7_4d29]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1345_c32_f967]
signal BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1345_c32_6bce]
signal BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1345_c32_bd93]
signal MUX_uxn_opcodes_h_l1345_c32_bd93_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1345_c32_bd93_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1345_c32_bd93_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1345_c32_bd93_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1347_c11_9000]
signal BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1347_c7_091d]
signal result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1347_c7_091d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1347_c7_091d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1347_c7_091d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1347_c7_091d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1351_c24_586d]
signal BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1353_c11_bf87]
signal BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1353_c7_d7a3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1353_c7_d7a3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_df93( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_value := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_stack_read := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_opc_done := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074
BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_left,
BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_right,
BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_return_output);

-- t8_MUX_uxn_opcodes_h_l1332_c2_0ed7
t8_MUX_uxn_opcodes_h_l1332_c2_0ed7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond,
t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue,
t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse,
t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7
result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond,
result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7
result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7
result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7
result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7
result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7
result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output);

-- printf_uxn_opcodes_h_l1333_c3_da23_uxn_opcodes_h_l1333_c3_da23
printf_uxn_opcodes_h_l1333_c3_da23_uxn_opcodes_h_l1333_c3_da23 : entity work.printf_uxn_opcodes_h_l1333_c3_da23_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1333_c3_da23_uxn_opcodes_h_l1333_c3_da23_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61
BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_left,
BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_right,
BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output);

-- t8_MUX_uxn_opcodes_h_l1338_c7_8e08
t8_MUX_uxn_opcodes_h_l1338_c7_8e08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1338_c7_8e08_cond,
t8_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue,
t8_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse,
t8_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08
result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_cond,
result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08
result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08
result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08
result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08
result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08
result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434
BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_left,
BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_right,
BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output);

-- t8_MUX_uxn_opcodes_h_l1341_c7_4d29
t8_MUX_uxn_opcodes_h_l1341_c7_4d29 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1341_c7_4d29_cond,
t8_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue,
t8_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse,
t8_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29
result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_cond,
result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29
result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29
result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29
result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29
result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29
result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967
BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_left,
BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_right,
BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce
BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_left,
BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_right,
BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_return_output);

-- MUX_uxn_opcodes_h_l1345_c32_bd93
MUX_uxn_opcodes_h_l1345_c32_bd93 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1345_c32_bd93_cond,
MUX_uxn_opcodes_h_l1345_c32_bd93_iftrue,
MUX_uxn_opcodes_h_l1345_c32_bd93_iffalse,
MUX_uxn_opcodes_h_l1345_c32_bd93_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000
BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_left,
BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_right,
BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d
result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_cond,
result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d
result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d
result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d
result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d
BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_left,
BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_right,
BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87
BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_left,
BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_right,
BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3
result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3
result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_return_output,
 t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output,
 t8_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output,
 t8_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_return_output,
 MUX_uxn_opcodes_h_l1345_c32_bd93_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1335_c3_b3f1 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1333_c3_da23_uxn_opcodes_h_l1333_c3_da23_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1339_c3_aa17 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1345_c32_bd93_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1345_c32_bd93_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1345_c32_bd93_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1345_c32_bd93_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_uxn_opcodes_h_l1351_c3_bdc3 : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1350_c3_0b41 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_return_output : unsigned(8 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1338_l1341_l1332_l1347_DUPLICATE_73b9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1338_l1332_l1347_DUPLICATE_7a67_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1338_l1341_l1332_DUPLICATE_8a66_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1332_DUPLICATE_2358_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1338_l1341_DUPLICATE_d9f8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1347_DUPLICATE_454e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1341_l1347_DUPLICATE_8cb1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_df93_uxn_opcodes_h_l1358_l1328_DUPLICATE_8c0c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_right := to_unsigned(0, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_right := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1345_c32_bd93_iffalse := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_right := to_unsigned(3, 2);
     VAR_BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_right := to_unsigned(2, 2);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_right := to_unsigned(128, 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1350_c3_0b41 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1350_c3_0b41;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1335_c3_b3f1 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1335_c3_b3f1;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1339_c3_aa17 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1339_c3_aa17;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1345_c32_bd93_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1338_l1341_l1332_l1347_DUPLICATE_73b9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1338_l1341_l1332_l1347_DUPLICATE_73b9_return_output := result.stack_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1332_c6_b074] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_left;
     BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output := BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1351_c24_586d] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1341_l1347_DUPLICATE_8cb1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1341_l1347_DUPLICATE_8cb1_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1338_l1341_l1332_DUPLICATE_8a66 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1338_l1341_l1332_DUPLICATE_8a66_return_output := result.sp_relative_shift;

     -- BIN_OP_AND[uxn_opcodes_h_l1345_c32_f967] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_left;
     BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_return_output := BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1353_c11_bf87] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_left;
     BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_return_output := BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1341_c11_0434] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_left;
     BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output := BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1338_l1332_l1347_DUPLICATE_7a67 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1338_l1332_l1347_DUPLICATE_7a67_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1338_l1341_DUPLICATE_d9f8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1338_l1341_DUPLICATE_d9f8_return_output := result.is_stack_read;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1347_DUPLICATE_454e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1347_DUPLICATE_454e_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1338_c11_3b61] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_left;
     BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output := BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1332_DUPLICATE_2358 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1332_DUPLICATE_2358_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1347_c11_9000] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_left;
     BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_return_output := BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1345_c32_f967_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c6_b074_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1338_c7_8e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c11_3b61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1341_c7_4d29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1341_c11_0434_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1347_c11_9000_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1353_c11_bf87_return_output;
     VAR_result_stack_value_uxn_opcodes_h_l1351_c3_bdc3 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1351_c24_586d_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1338_l1341_l1332_DUPLICATE_8a66_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1338_l1341_l1332_DUPLICATE_8a66_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1338_l1341_l1332_DUPLICATE_8a66_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1347_DUPLICATE_454e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1347_DUPLICATE_454e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1347_DUPLICATE_454e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1347_DUPLICATE_454e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1338_l1332_l1347_DUPLICATE_7a67_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1338_l1332_l1347_DUPLICATE_7a67_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1338_l1332_l1347_DUPLICATE_7a67_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1338_l1341_DUPLICATE_d9f8_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1338_l1341_DUPLICATE_d9f8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1332_DUPLICATE_2358_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1332_DUPLICATE_2358_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1332_DUPLICATE_2358_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1338_l1353_l1341_l1332_DUPLICATE_2358_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1341_l1347_DUPLICATE_8cb1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1341_l1347_DUPLICATE_8cb1_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1338_l1341_l1332_l1347_DUPLICATE_73b9_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1338_l1341_l1332_l1347_DUPLICATE_73b9_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1338_l1341_l1332_l1347_DUPLICATE_73b9_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1338_l1341_l1332_l1347_DUPLICATE_73b9_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue := VAR_result_stack_value_uxn_opcodes_h_l1351_c3_bdc3;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1353_c7_d7a3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1353_c7_d7a3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1347_c7_091d] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_return_output := result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1347_c7_091d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1332_c1_5c08] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1347_c7_091d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_return_output;

     -- t8_MUX[uxn_opcodes_h_l1341_c7_4d29] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1341_c7_4d29_cond <= VAR_t8_MUX_uxn_opcodes_h_l1341_c7_4d29_cond;
     t8_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue;
     t8_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output := t8_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1341_c7_4d29] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1345_c32_6bce] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_left;
     BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_return_output := BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1345_c32_bd93_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1345_c32_6bce_return_output;
     VAR_printf_uxn_opcodes_h_l1333_c3_da23_uxn_opcodes_h_l1333_c3_da23_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1332_c1_5c08_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1347_c7_091d_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1353_c7_d7a3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1347_c7_091d_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1347_c7_091d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;
     -- printf_uxn_opcodes_h_l1333_c3_da23[uxn_opcodes_h_l1333_c3_da23] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1333_c3_da23_uxn_opcodes_h_l1333_c3_da23_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1333_c3_da23_uxn_opcodes_h_l1333_c3_da23_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1347_c7_091d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_return_output;

     -- MUX[uxn_opcodes_h_l1345_c32_bd93] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1345_c32_bd93_cond <= VAR_MUX_uxn_opcodes_h_l1345_c32_bd93_cond;
     MUX_uxn_opcodes_h_l1345_c32_bd93_iftrue <= VAR_MUX_uxn_opcodes_h_l1345_c32_bd93_iftrue;
     MUX_uxn_opcodes_h_l1345_c32_bd93_iffalse <= VAR_MUX_uxn_opcodes_h_l1345_c32_bd93_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1345_c32_bd93_return_output := MUX_uxn_opcodes_h_l1345_c32_bd93_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1341_c7_4d29] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1338_c7_8e08] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1347_c7_091d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_return_output;

     -- t8_MUX[uxn_opcodes_h_l1338_c7_8e08] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1338_c7_8e08_cond <= VAR_t8_MUX_uxn_opcodes_h_l1338_c7_8e08_cond;
     t8_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue;
     t8_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output := t8_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1341_c7_4d29] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1341_c7_4d29] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output := result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue := VAR_MUX_uxn_opcodes_h_l1345_c32_bd93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1347_c7_091d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1347_c7_091d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1338_c7_8e08] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;

     -- t8_MUX[uxn_opcodes_h_l1332_c2_0ed7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond <= VAR_t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond;
     t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue;
     t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output := t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1341_c7_4d29] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1338_c7_8e08] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1332_c2_0ed7] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1341_c7_4d29] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1338_c7_8e08] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output := result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1341_c7_4d29] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1341_c7_4d29_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1338_c7_8e08] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1332_c2_0ed7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1332_c2_0ed7] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output := result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1338_c7_8e08] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1338_c7_8e08] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1332_c2_0ed7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1338_c7_8e08_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1332_c2_0ed7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1332_c2_0ed7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1332_c2_0ed7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_df93_uxn_opcodes_h_l1358_l1328_DUPLICATE_8c0c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_df93_uxn_opcodes_h_l1358_l1328_DUPLICATE_8c0c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_df93(
     result,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c2_0ed7_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_df93_uxn_opcodes_h_l1358_l1328_DUPLICATE_8c0c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_df93_uxn_opcodes_h_l1358_l1328_DUPLICATE_8c0c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
