-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity equ_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_226c8821;
architecture arch of equ_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1162_c6_4531]
signal BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1162_c2_6c56]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1162_c2_6c56]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1162_c2_6c56]
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1162_c2_6c56]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1162_c2_6c56]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1162_c2_6c56]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1162_c2_6c56]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1162_c2_6c56]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1162_c2_6c56]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1162_c2_6c56]
signal n8_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1162_c2_6c56]
signal t8_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1175_c11_2d93]
signal BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1175_c7_de44]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1175_c7_de44]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1175_c7_de44]
signal result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1175_c7_de44]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1175_c7_de44]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1175_c7_de44]
signal n8_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1175_c7_de44]
signal t8_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1178_c11_6c24]
signal BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1178_c7_5387]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1178_c7_5387]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1178_c7_5387]
signal result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1178_c7_5387]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1178_c7_5387]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1178_c7_5387]
signal n8_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1178_c7_5387]
signal t8_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1181_c11_38f3]
signal BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1181_c7_824c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1181_c7_824c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1181_c7_824c]
signal result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1181_c7_824c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1181_c7_824c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1181_c7_824c]
signal n8_MUX_uxn_opcodes_h_l1181_c7_824c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1181_c7_824c_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1183_c30_1c08]
signal sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1186_c21_a8b9]
signal BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1186_c21_9ea5]
signal MUX_uxn_opcodes_h_l1186_c21_9ea5_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1186_c21_9ea5_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1186_c21_9ea5_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1186_c21_9ea5_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_left,
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_right,
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_cond,
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output);

-- n8_MUX_uxn_opcodes_h_l1162_c2_6c56
n8_MUX_uxn_opcodes_h_l1162_c2_6c56 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1162_c2_6c56_cond,
n8_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue,
n8_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse,
n8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output);

-- t8_MUX_uxn_opcodes_h_l1162_c2_6c56
t8_MUX_uxn_opcodes_h_l1162_c2_6c56 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1162_c2_6c56_cond,
t8_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue,
t8_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse,
t8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93
BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_left,
BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_right,
BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_cond,
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_return_output);

-- n8_MUX_uxn_opcodes_h_l1175_c7_de44
n8_MUX_uxn_opcodes_h_l1175_c7_de44 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1175_c7_de44_cond,
n8_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue,
n8_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse,
n8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output);

-- t8_MUX_uxn_opcodes_h_l1175_c7_de44
t8_MUX_uxn_opcodes_h_l1175_c7_de44 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1175_c7_de44_cond,
t8_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue,
t8_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse,
t8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24
BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_left,
BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_right,
BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_cond,
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_return_output);

-- n8_MUX_uxn_opcodes_h_l1178_c7_5387
n8_MUX_uxn_opcodes_h_l1178_c7_5387 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1178_c7_5387_cond,
n8_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue,
n8_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse,
n8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output);

-- t8_MUX_uxn_opcodes_h_l1178_c7_5387
t8_MUX_uxn_opcodes_h_l1178_c7_5387 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1178_c7_5387_cond,
t8_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue,
t8_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse,
t8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3
BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_left,
BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_right,
BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_return_output);

-- n8_MUX_uxn_opcodes_h_l1181_c7_824c
n8_MUX_uxn_opcodes_h_l1181_c7_824c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1181_c7_824c_cond,
n8_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue,
n8_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse,
n8_MUX_uxn_opcodes_h_l1181_c7_824c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08
sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_ins,
sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_x,
sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_y,
sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9
BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_left,
BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_right,
BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_return_output);

-- MUX_uxn_opcodes_h_l1186_c21_9ea5
MUX_uxn_opcodes_h_l1186_c21_9ea5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1186_c21_9ea5_cond,
MUX_uxn_opcodes_h_l1186_c21_9ea5_iftrue,
MUX_uxn_opcodes_h_l1186_c21_9ea5_iffalse,
MUX_uxn_opcodes_h_l1186_c21_9ea5_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
 n8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
 t8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_return_output,
 n8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output,
 t8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_return_output,
 n8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output,
 t8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_return_output,
 n8_MUX_uxn_opcodes_h_l1181_c7_824c_return_output,
 sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_return_output,
 MUX_uxn_opcodes_h_l1186_c21_9ea5_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1167_c3_1a08 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1172_c3_ccc3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1162_c2_6c56_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1176_c3_a47f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1175_c7_de44_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1181_c7_824c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5387_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1185_c3_4f09 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1181_c7_824c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1186_c21_9ea5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1186_c21_9ea5_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1186_c21_9ea5_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1186_c21_9ea5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1178_l1162_l1181_l1175_DUPLICATE_3a06_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_40cd_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_f377_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_286e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1178_l1181_DUPLICATE_bb79_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1190_l1158_DUPLICATE_ee9a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1176_c3_a47f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1176_c3_a47f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1172_c3_ccc3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1172_c3_ccc3;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1186_c21_9ea5_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1185_c3_4f09 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1185_c3_4f09;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1167_c3_1a08 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1167_c3_1a08;
     VAR_MUX_uxn_opcodes_h_l1186_c21_9ea5_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1175_c11_2d93] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_left;
     BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_return_output := BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1181_c11_38f3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1162_c2_6c56_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1162_c6_4531] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_left;
     BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output := BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1178_l1162_l1181_l1175_DUPLICATE_3a06 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1178_l1162_l1181_l1175_DUPLICATE_3a06_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1186_c21_a8b9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1178_l1181_DUPLICATE_bb79 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1178_l1181_DUPLICATE_bb79_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1162_c2_6c56_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_f377 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_f377_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1178_c11_6c24] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_left;
     BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_return_output := BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1183_c30_1c08] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_ins;
     sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_x;
     sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_return_output := sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1162_c2_6c56_return_output := result.is_vram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_40cd LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_40cd_return_output := result.sp_relative_shift;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1162_c2_6c56_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_286e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_286e_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1162_c2_6c56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1162_c2_6c56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_4531_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1175_c7_de44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1175_c7_de44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1175_c11_2d93_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1178_c11_6c24_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1181_c7_824c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1181_c11_38f3_return_output;
     VAR_MUX_uxn_opcodes_h_l1186_c21_9ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c21_a8b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_40cd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_40cd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_40cd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_286e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_286e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_286e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_f377_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_f377_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1178_l1181_l1175_DUPLICATE_f377_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1178_l1181_DUPLICATE_bb79_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1178_l1181_DUPLICATE_bb79_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1178_l1162_l1181_l1175_DUPLICATE_3a06_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1178_l1162_l1181_l1175_DUPLICATE_3a06_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1178_l1162_l1181_l1175_DUPLICATE_3a06_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1178_l1162_l1181_l1175_DUPLICATE_3a06_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1162_c2_6c56_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1162_c2_6c56_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1162_c2_6c56_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1162_c2_6c56_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1183_c30_1c08_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output;

     -- n8_MUX[uxn_opcodes_h_l1181_c7_824c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1181_c7_824c_cond <= VAR_n8_MUX_uxn_opcodes_h_l1181_c7_824c_cond;
     n8_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue;
     n8_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1181_c7_824c_return_output := n8_MUX_uxn_opcodes_h_l1181_c7_824c_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1181_c7_824c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1181_c7_824c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1181_c7_824c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1178_c7_5387] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1178_c7_5387_cond <= VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5387_cond;
     t8_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue;
     t8_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output := t8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1181_c7_824c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output;

     -- MUX[uxn_opcodes_h_l1186_c21_9ea5] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1186_c21_9ea5_cond <= VAR_MUX_uxn_opcodes_h_l1186_c21_9ea5_cond;
     MUX_uxn_opcodes_h_l1186_c21_9ea5_iftrue <= VAR_MUX_uxn_opcodes_h_l1186_c21_9ea5_iftrue;
     MUX_uxn_opcodes_h_l1186_c21_9ea5_iffalse <= VAR_MUX_uxn_opcodes_h_l1186_c21_9ea5_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1186_c21_9ea5_return_output := MUX_uxn_opcodes_h_l1186_c21_9ea5_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue := VAR_MUX_uxn_opcodes_h_l1186_c21_9ea5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1181_c7_824c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1181_c7_824c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1181_c7_824c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1181_c7_824c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1181_c7_824c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;
     -- n8_MUX[uxn_opcodes_h_l1178_c7_5387] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1178_c7_5387_cond <= VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5387_cond;
     n8_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue;
     n8_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output := n8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1181_c7_824c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1178_c7_5387] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1178_c7_5387] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;

     -- t8_MUX[uxn_opcodes_h_l1175_c7_de44] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1175_c7_de44_cond <= VAR_t8_MUX_uxn_opcodes_h_l1175_c7_de44_cond;
     t8_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue;
     t8_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output := t8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1178_c7_5387] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1178_c7_5387] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1181_c7_824c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1175_c7_de44] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1178_c7_5387] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_return_output := result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;

     -- t8_MUX[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1162_c2_6c56_cond <= VAR_t8_MUX_uxn_opcodes_h_l1162_c2_6c56_cond;
     t8_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue;
     t8_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output := t8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1175_c7_de44] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;

     -- n8_MUX[uxn_opcodes_h_l1175_c7_de44] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1175_c7_de44_cond <= VAR_n8_MUX_uxn_opcodes_h_l1175_c7_de44_cond;
     n8_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue;
     n8_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output := n8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1175_c7_de44] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1175_c7_de44] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1178_c7_5387_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output;

     -- n8_MUX[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1162_c2_6c56_cond <= VAR_n8_MUX_uxn_opcodes_h_l1162_c2_6c56_cond;
     n8_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue;
     n8_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output := n8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1175_c7_de44] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_return_output := result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1175_c7_de44_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1162_c2_6c56] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output := result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1190_l1158_DUPLICATE_ee9a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1190_l1158_DUPLICATE_ee9a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_6c56_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1190_l1158_DUPLICATE_ee9a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1190_l1158_DUPLICATE_ee9a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
