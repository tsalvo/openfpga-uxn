-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity rot_0CLK_af0b7c12 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end rot_0CLK_af0b7c12;
architecture arch of rot_0CLK_af0b7c12 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2361_c6_dad8]
signal BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2361_c2_1656]
signal l8_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2361_c2_1656]
signal result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2361_c2_1656]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2361_c2_1656]
signal result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2361_c2_1656]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2361_c2_1656]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2361_c2_1656]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2361_c2_1656]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2361_c2_1656]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2361_c2_1656]
signal tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2369_c11_4af8]
signal BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2369_c7_eafd]
signal l8_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2369_c7_eafd]
signal result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2369_c7_eafd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2369_c7_eafd]
signal result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2369_c7_eafd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2369_c7_eafd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2369_c7_eafd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2369_c7_eafd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2369_c7_eafd]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2369_c7_eafd]
signal tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2373_c11_e7ff]
signal BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2373_c7_2f7e]
signal l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2373_c7_2f7e]
signal result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2373_c7_2f7e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2373_c7_2f7e]
signal result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2373_c7_2f7e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2373_c7_2f7e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2373_c7_2f7e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2373_c7_2f7e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2373_c7_2f7e]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l2373_c7_2f7e]
signal tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2376_c30_d3ae]
signal sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2382_c11_d5d4]
signal BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2382_c7_46d5]
signal l8_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2382_c7_46d5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2382_c7_46d5]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2382_c7_46d5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2382_c7_46d5]
signal result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2382_c7_46d5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2382_c7_46d5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2389_c11_e99e]
signal BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2389_c7_fedd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2389_c7_fedd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_4982( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_sp_shift := ref_toks_7;
      base.is_stack_operation_16bit := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8
BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_left,
BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_right,
BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output);

-- l8_MUX_uxn_opcodes_h_l2361_c2_1656
l8_MUX_uxn_opcodes_h_l2361_c2_1656 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2361_c2_1656_cond,
l8_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue,
l8_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse,
l8_MUX_uxn_opcodes_h_l2361_c2_1656_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656
result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_cond,
result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656
result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656
result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_cond,
result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656
result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656
result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656
result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2361_c2_1656
tmp16_MUX_uxn_opcodes_h_l2361_c2_1656 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_cond,
tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue,
tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse,
tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8
BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_left,
BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_right,
BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output);

-- l8_MUX_uxn_opcodes_h_l2369_c7_eafd
l8_MUX_uxn_opcodes_h_l2369_c7_eafd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2369_c7_eafd_cond,
l8_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue,
l8_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse,
l8_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd
result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_cond,
result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd
result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd
result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_cond,
result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd
result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd
result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd
result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd
tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_cond,
tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue,
tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse,
tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff
BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_left,
BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_right,
BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output);

-- l8_MUX_uxn_opcodes_h_l2373_c7_2f7e
l8_MUX_uxn_opcodes_h_l2373_c7_2f7e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond,
l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue,
l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse,
l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e
result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond,
result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e
result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e
result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e
result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e
result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output);

-- tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e
tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond,
tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue,
tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse,
tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae
sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_ins,
sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_x,
sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_y,
sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4
BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_left,
BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_right,
BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_return_output);

-- l8_MUX_uxn_opcodes_h_l2382_c7_46d5
l8_MUX_uxn_opcodes_h_l2382_c7_46d5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2382_c7_46d5_cond,
l8_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue,
l8_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse,
l8_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5
result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5
result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5
result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_cond,
result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5
result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e
BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_left,
BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_right,
BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd
result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd
result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 tmp16,
 t8,
 n8,
 l8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output,
 l8_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
 tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output,
 l8_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output,
 tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output,
 l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output,
 tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output,
 sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_return_output,
 l8_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2366_c3_1f12 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2370_c3_2857 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2379_c3_a659 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2386_c3_a70e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2382_c7_46d5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2383_c8_a94b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2373_l2361_l2369_DUPLICATE_ee6c_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2373_l2361_l2382_l2369_DUPLICATE_dd4d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2373_l2361_l2369_DUPLICATE_a4ec_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2361_l2382_l2369_l2389_DUPLICATE_55d6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2361_l2382_l2369_DUPLICATE_2127_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2373_l2382_l2369_l2389_DUPLICATE_4e44_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4982_uxn_opcodes_h_l2394_l2356_DUPLICATE_35ff_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_tmp16 := tmp16;
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2366_c3_1f12 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2366_c3_1f12;
     VAR_sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2370_c3_2857 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2370_c3_2857;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2379_c3_a659 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2379_c3_a659;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2386_c3_a70e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2386_c3_a70e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_right := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_ins := VAR_ins;
     VAR_l8_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse := l8;
     REG_VAR_n8 := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_left := VAR_phase;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue := VAR_previous_stack_read;
     VAR_tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue := VAR_previous_stack_read;
     REG_VAR_t8 := t8;
     VAR_tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse := tmp16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2361_l2382_l2369_DUPLICATE_2127 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2361_l2382_l2369_DUPLICATE_2127_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2373_c11_e7ff] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_left;
     BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output := BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2382_c7_46d5] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2382_c7_46d5_return_output := result.stack_address_sp_offset;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2383_c8_a94b] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2383_c8_a94b_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l2369_c11_4af8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2382_c11_d5d4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2361_l2382_l2369_l2389_DUPLICATE_55d6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2361_l2382_l2369_l2389_DUPLICATE_55d6_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2389_c11_e99e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_return_output;

     -- result_is_stack_operation_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d[uxn_opcodes_h_l2382_c7_46d5] LATENCY=0
     VAR_result_is_stack_operation_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2382_c7_46d5_return_output := result.is_stack_operation_16bit;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2373_l2382_l2369_l2389_DUPLICATE_4e44 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2373_l2382_l2369_l2389_DUPLICATE_4e44_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2373_l2361_l2369_DUPLICATE_ee6c LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2373_l2361_l2369_DUPLICATE_ee6c_return_output := result.u16_value;

     -- sp_relative_shift[uxn_opcodes_h_l2376_c30_d3ae] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_ins;
     sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_x;
     sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_return_output := sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2373_l2361_l2382_l2369_DUPLICATE_dd4d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2373_l2361_l2382_l2369_DUPLICATE_dd4d_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2361_c6_dad8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2373_l2361_l2369_DUPLICATE_a4ec LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2373_l2361_l2369_DUPLICATE_a4ec_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_l8_MUX_uxn_opcodes_h_l2361_c2_1656_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2361_c6_dad8_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2369_c7_eafd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2369_c11_4af8_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2373_c11_e7ff_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2382_c7_46d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2382_c11_d5d4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2389_c11_e99e_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2383_c8_a94b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2383_c8_a94b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2373_l2361_l2369_DUPLICATE_a4ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2373_l2361_l2369_DUPLICATE_a4ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2373_l2361_l2369_DUPLICATE_a4ec_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2373_l2361_l2369_DUPLICATE_ee6c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2373_l2361_l2369_DUPLICATE_ee6c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2373_l2361_l2369_DUPLICATE_ee6c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2373_l2382_l2369_l2389_DUPLICATE_4e44_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2373_l2382_l2369_l2389_DUPLICATE_4e44_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2373_l2382_l2369_l2389_DUPLICATE_4e44_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2373_l2382_l2369_l2389_DUPLICATE_4e44_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2361_l2382_l2369_DUPLICATE_2127_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2361_l2382_l2369_DUPLICATE_2127_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2361_l2382_l2369_DUPLICATE_2127_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2361_l2382_l2369_l2389_DUPLICATE_55d6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2361_l2382_l2369_l2389_DUPLICATE_55d6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2361_l2382_l2369_l2389_DUPLICATE_55d6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2361_l2382_l2369_l2389_DUPLICATE_55d6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2373_l2361_l2382_l2369_DUPLICATE_dd4d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2373_l2361_l2382_l2369_DUPLICATE_dd4d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2373_l2361_l2382_l2369_DUPLICATE_dd4d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2373_l2361_l2382_l2369_DUPLICATE_dd4d_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse := VAR_result_is_stack_operation_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2382_c7_46d5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2382_c7_46d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2376_c30_d3ae_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2373_c7_2f7e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2382_c7_46d5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output := result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2382_c7_46d5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2382_c7_46d5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;

     -- l8_MUX[uxn_opcodes_h_l2382_c7_46d5] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2382_c7_46d5_cond <= VAR_l8_MUX_uxn_opcodes_h_l2382_c7_46d5_cond;
     l8_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue;
     l8_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output := l8_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l2373_c7_2f7e] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond;
     tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output := tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2382_c7_46d5] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2389_c7_fedd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2373_c7_2f7e] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output := result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2389_c7_fedd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output;

     -- Submodule level 2
     VAR_l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2389_c7_fedd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2373_c7_2f7e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2369_c7_eafd] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output := result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l2369_c7_eafd] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_cond;
     tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output := tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2382_c7_46d5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2373_c7_2f7e] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;

     -- l8_MUX[uxn_opcodes_h_l2373_c7_2f7e] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond <= VAR_l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond;
     l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue;
     l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output := l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2369_c7_eafd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2373_c7_2f7e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2373_c7_2f7e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2382_c7_46d5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;

     -- Submodule level 3
     VAR_l8_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2382_c7_46d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2373_c7_2f7e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2369_c7_eafd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2369_c7_eafd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output := result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2361_c2_1656] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2369_c7_eafd] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2369_c7_eafd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2373_c7_2f7e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l2361_c2_1656] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_cond;
     tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue;
     tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_return_output := tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2361_c2_1656] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output := result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output;

     -- l8_MUX[uxn_opcodes_h_l2369_c7_eafd] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2369_c7_eafd_cond <= VAR_l8_MUX_uxn_opcodes_h_l2369_c7_eafd_cond;
     l8_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue;
     l8_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output := l8_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;

     -- Submodule level 4
     VAR_l8_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2373_c7_2f7e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l2361_c2_1656_return_output;
     -- l8_MUX[uxn_opcodes_h_l2361_c2_1656] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2361_c2_1656_cond <= VAR_l8_MUX_uxn_opcodes_h_l2361_c2_1656_cond;
     l8_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue;
     l8_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2361_c2_1656_return_output := l8_MUX_uxn_opcodes_h_l2361_c2_1656_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2369_c7_eafd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2361_c2_1656] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output := result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2361_c2_1656] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2361_c2_1656] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2369_c7_eafd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2361_c2_1656] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output;

     -- Submodule level 5
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l2361_c2_1656_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2369_c7_eafd_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2361_c2_1656] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2361_c2_1656] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4982_uxn_opcodes_h_l2394_l2356_DUPLICATE_35ff LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4982_uxn_opcodes_h_l2394_l2356_DUPLICATE_35ff_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4982(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2361_c2_1656_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2361_c2_1656_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4982_uxn_opcodes_h_l2394_l2356_DUPLICATE_35ff_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4982_uxn_opcodes_h_l2394_l2356_DUPLICATE_35ff_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     tmp16 <= REG_COMB_tmp16;
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
