-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 35
entity dup_0CLK_02ab8d09 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_02ab8d09;
architecture arch of dup_0CLK_02ab8d09 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2956_c6_f36b]
signal BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2956_c2_0c8c]
signal t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2956_c2_0c8c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2956_c2_0c8c]
signal result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2956_c2_0c8c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2956_c2_0c8c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2956_c2_0c8c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2956_c2_0c8c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2961_c11_39e8]
signal BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2961_c7_a8b3]
signal t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2961_c7_a8b3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2961_c7_a8b3]
signal result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2961_c7_a8b3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2961_c7_a8b3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2961_c7_a8b3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2961_c7_a8b3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2964_c11_e352]
signal BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2964_c7_dc8a]
signal t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2964_c7_dc8a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2964_c7_dc8a]
signal result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2964_c7_dc8a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2964_c7_dc8a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2964_c7_dc8a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2964_c7_dc8a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2967_c30_611b]
signal sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2972_c11_4b8b]
signal BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2972_c7_af11]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2972_c7_af11]
signal result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2972_c7_af11]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2972_c7_af11]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2972_c7_af11]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2977_c11_4154]
signal BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2977_c7_767f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2977_c7_767f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_3345( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b
BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_left,
BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_right,
BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_return_output);

-- t8_MUX_uxn_opcodes_h_l2956_c2_0c8c
t8_MUX_uxn_opcodes_h_l2956_c2_0c8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond,
t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue,
t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse,
t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c
result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c
result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c
result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c
result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8
BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_left,
BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_right,
BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_return_output);

-- t8_MUX_uxn_opcodes_h_l2961_c7_a8b3
t8_MUX_uxn_opcodes_h_l2961_c7_a8b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond,
t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue,
t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse,
t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3
result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3
result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3
result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3
result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352
BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_left,
BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_right,
BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_return_output);

-- t8_MUX_uxn_opcodes_h_l2964_c7_dc8a
t8_MUX_uxn_opcodes_h_l2964_c7_dc8a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond,
t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue,
t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse,
t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a
result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a
result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a
result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a
result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2967_c30_611b
sp_relative_shift_uxn_opcodes_h_l2967_c30_611b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_ins,
sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_x,
sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_y,
sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b
BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_left,
BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_right,
BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11
result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_cond,
result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11
result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11
result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11
result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154
BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_left,
BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_right,
BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f
result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f
result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_return_output,
 t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_return_output,
 t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_return_output,
 t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output,
 sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2958_c3_385a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2962_c3_2fde : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2969_c3_31bc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2974_c3_a5bd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2972_c7_af11_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2961_l2956_l2972_DUPLICATE_d238_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2961_l2977_l2956_l2972_DUPLICATE_d2b2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2961_l2964_l2956_DUPLICATE_8828_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2961_l2956_l2972_DUPLICATE_811e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2977_l2964_l2972_DUPLICATE_4a87_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2952_l2982_DUPLICATE_fe8a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2969_c3_31bc := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2969_c3_31bc;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2962_c3_2fde := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2962_c3_2fde;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2958_c3_385a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2958_c3_385a;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2974_c3_a5bd := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2974_c3_a5bd;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2961_l2964_l2956_DUPLICATE_8828 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2961_l2964_l2956_DUPLICATE_8828_return_output := result.sp_relative_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2972_c7_af11] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2972_c7_af11_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2977_c11_4154] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_left;
     BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_return_output := BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2956_c6_f36b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2961_c11_39e8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2972_c11_4b8b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2964_c11_e352] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_left;
     BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_return_output := BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2961_l2956_l2972_DUPLICATE_811e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2961_l2956_l2972_DUPLICATE_811e_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2961_l2956_l2972_DUPLICATE_d238 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2961_l2956_l2972_DUPLICATE_d238_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2961_l2977_l2956_l2972_DUPLICATE_d2b2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2961_l2977_l2956_l2972_DUPLICATE_d2b2_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l2967_c30_611b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_ins;
     sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_x;
     sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_return_output := sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2977_l2964_l2972_DUPLICATE_4a87 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2977_l2964_l2972_DUPLICATE_4a87_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2956_c6_f36b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_39e8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2964_c11_e352_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2972_c11_4b8b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2977_c11_4154_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2961_l2964_l2956_DUPLICATE_8828_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2961_l2964_l2956_DUPLICATE_8828_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2961_l2964_l2956_DUPLICATE_8828_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2977_l2964_l2972_DUPLICATE_4a87_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2977_l2964_l2972_DUPLICATE_4a87_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2977_l2964_l2972_DUPLICATE_4a87_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2977_l2964_l2972_DUPLICATE_4a87_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2961_l2956_l2972_DUPLICATE_811e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2961_l2956_l2972_DUPLICATE_811e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2961_l2956_l2972_DUPLICATE_811e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2961_l2977_l2956_l2972_DUPLICATE_d2b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2961_l2977_l2956_l2972_DUPLICATE_d2b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2961_l2977_l2956_l2972_DUPLICATE_d2b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2961_l2977_l2956_l2972_DUPLICATE_d2b2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2961_l2956_l2972_DUPLICATE_d238_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2961_l2956_l2972_DUPLICATE_d238_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2961_l2956_l2972_DUPLICATE_d238_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2972_c7_af11_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2967_c30_611b_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2972_c7_af11] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2977_c7_767f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2964_c7_dc8a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2977_c7_767f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2972_c7_af11] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_return_output := result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_return_output;

     -- t8_MUX[uxn_opcodes_h_l2964_c7_dc8a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond <= VAR_t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond;
     t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue;
     t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output := t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2972_c7_af11] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2977_c7_767f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2972_c7_af11_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2977_c7_767f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2972_c7_af11_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2972_c7_af11_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2961_c7_a8b3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2964_c7_dc8a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;

     -- t8_MUX[uxn_opcodes_h_l2961_c7_a8b3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond <= VAR_t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond;
     t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue;
     t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output := t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2964_c7_dc8a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2964_c7_dc8a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2972_c7_af11] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2972_c7_af11] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2972_c7_af11_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2972_c7_af11_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2964_c7_dc8a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2956_c2_0c8c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2961_c7_a8b3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2961_c7_a8b3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2964_c7_dc8a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2961_c7_a8b3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;

     -- t8_MUX[uxn_opcodes_h_l2956_c2_0c8c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond <= VAR_t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond;
     t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue;
     t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output := t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2964_c7_dc8a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2961_c7_a8b3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2961_c7_a8b3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2956_c2_0c8c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2956_c2_0c8c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2956_c2_0c8c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_a8b3_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2956_c2_0c8c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2956_c2_0c8c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2952_l2982_DUPLICATE_fe8a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2952_l2982_DUPLICATE_fe8a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3345(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2956_c2_0c8c_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2952_l2982_DUPLICATE_fe8a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2952_l2982_DUPLICATE_fe8a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
