-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 11
entity opc_pop2_phased_0CLK_ba40181c is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_pop2_phased_0CLK_ba40181c;
architecture arch of opc_pop2_phased_0CLK_ba40181c is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal set_will_succeed : unsigned(0 downto 0) := to_unsigned(0, 1);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_set_will_succeed : unsigned(0 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l193_c6_cd6a]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l193_c1_c261]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l196_c7_11a1]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l193_c2_d23e]
signal result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_return_output : unsigned(0 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l194_c12_f63a]
signal set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l196_c11_85bd]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l196_c1_8293]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l196_c7_11a1]
signal result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output : unsigned(0 downto 0);

-- set[uxn_opcodes_phased_h_l197_c3_b6cd]
signal set_uxn_opcodes_phased_h_l197_c3_b6cd_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l197_c3_b6cd_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l197_c3_b6cd_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l197_c3_b6cd_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l197_c3_b6cd_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l197_c3_b6cd_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l197_c3_b6cd_add : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l199_c11_a415]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l199_c7_4894]
signal result_MUX_uxn_opcodes_phased_h_l199_c7_4894_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l199_c7_4894_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l199_c7_4894_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l199_c7_4894_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a
BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output);

-- result_MUX_uxn_opcodes_phased_h_l193_c2_d23e
result_MUX_uxn_opcodes_phased_h_l193_c2_d23e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_cond,
result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_iftrue,
result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_iffalse,
result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a
set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_sp,
set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_k,
set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_mul,
set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_add,
set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd
BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_return_output);

-- result_MUX_uxn_opcodes_phased_h_l196_c7_11a1
result_MUX_uxn_opcodes_phased_h_l196_c7_11a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_cond,
result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iftrue,
result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iffalse,
result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output);

-- set_uxn_opcodes_phased_h_l197_c3_b6cd
set_uxn_opcodes_phased_h_l197_c3_b6cd : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l197_c3_b6cd_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l197_c3_b6cd_sp,
set_uxn_opcodes_phased_h_l197_c3_b6cd_stack_index,
set_uxn_opcodes_phased_h_l197_c3_b6cd_ins,
set_uxn_opcodes_phased_h_l197_c3_b6cd_k,
set_uxn_opcodes_phased_h_l197_c3_b6cd_mul,
set_uxn_opcodes_phased_h_l197_c3_b6cd_add);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415
BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_return_output);

-- result_MUX_uxn_opcodes_phased_h_l199_c7_4894
result_MUX_uxn_opcodes_phased_h_l199_c7_4894 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l199_c7_4894_cond,
result_MUX_uxn_opcodes_phased_h_l199_c7_4894_iftrue,
result_MUX_uxn_opcodes_phased_h_l199_c7_4894_iffalse,
result_MUX_uxn_opcodes_phased_h_l199_c7_4894_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 set_will_succeed,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output,
 result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_return_output,
 set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_return_output,
 result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_return_output,
 result_MUX_uxn_opcodes_phased_h_l199_c7_4894_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l199_c7_4894_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_cond : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l199_c7_4894_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l199_c7_4894_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l199_c7_4894_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_set_will_succeed : unsigned(0 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_set_will_succeed := set_will_succeed;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_MUX_uxn_opcodes_phased_h_l199_c7_4894_iftrue := to_unsigned(1, 1);
     VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_add := resize(to_signed(-2, 3), 8);
     VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_mul := resize(to_unsigned(2, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_right := to_unsigned(2, 2);
     VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_mul := resize(to_unsigned(2, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_iffalse := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_add := resize(to_signed(-2, 3), 8);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_k := VAR_k;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_left := VAR_phase;
     VAR_result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l199_c7_4894_iffalse := result;
     REG_VAR_set_will_succeed := set_will_succeed;
     VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_sp := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_stack_index := VAR_stack_index;
     -- BIN_OP_EQ[uxn_opcodes_phased_h_l196_c11_85bd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l193_c6_cd6a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l199_c11_a415] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l193_c6_cd6a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l196_c11_85bd_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l199_c7_4894_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l199_c11_a415_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l193_c1_c261] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l196_c7_11a1] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l199_c7_4894] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l199_c7_4894_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l199_c7_4894_cond;
     result_MUX_uxn_opcodes_phased_h_l199_c7_4894_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l199_c7_4894_iftrue;
     result_MUX_uxn_opcodes_phased_h_l199_c7_4894_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l199_c7_4894_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l199_c7_4894_return_output := result_MUX_uxn_opcodes_phased_h_l199_c7_4894_return_output;

     -- Submodule level 2
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l193_c1_c261_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l199_c7_4894_return_output;
     -- set_will_fail[uxn_opcodes_phased_h_l194_c12_f63a] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_sp;
     set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_k;
     set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_mul;
     set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_return_output := set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l196_c1_8293] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l196_c7_11a1] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_cond;
     result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iftrue;
     result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output := result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output;

     -- Submodule level 3
     VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l196_c1_8293_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l196_c7_11a1_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l194_c12_f63a_return_output;
     -- set[uxn_opcodes_phased_h_l197_c3_b6cd] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l197_c3_b6cd_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l197_c3_b6cd_sp <= VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_sp;
     set_uxn_opcodes_phased_h_l197_c3_b6cd_stack_index <= VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_stack_index;
     set_uxn_opcodes_phased_h_l197_c3_b6cd_ins <= VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_ins;
     set_uxn_opcodes_phased_h_l197_c3_b6cd_k <= VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_k;
     set_uxn_opcodes_phased_h_l197_c3_b6cd_mul <= VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_mul;
     set_uxn_opcodes_phased_h_l197_c3_b6cd_add <= VAR_set_uxn_opcodes_phased_h_l197_c3_b6cd_add;
     -- Outputs

     -- result_MUX[uxn_opcodes_phased_h_l193_c2_d23e] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_cond;
     result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_iftrue;
     result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_return_output := result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_return_output;

     -- Submodule level 4
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l193_c2_d23e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_set_will_succeed <= REG_VAR_set_will_succeed;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     set_will_succeed <= REG_COMB_set_will_succeed;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
