-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 54
entity div_0CLK_af9273cc is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end div_0CLK_af9273cc;
architecture arch of div_0CLK_af9273cc is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2190_c6_bf77]
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2190_c1_9bdd]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c2_91ed]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2190_c2_91ed]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c2_91ed]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c2_91ed]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2190_c2_91ed]
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c2_91ed]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2190_c2_91ed]
signal t8_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2190_c2_91ed]
signal n8_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2191_c3_4034[uxn_opcodes_h_l2191_c3_4034]
signal printf_uxn_opcodes_h_l2191_c3_4034_uxn_opcodes_h_l2191_c3_4034_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2195_c11_15a5]
signal BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2195_c7_45c6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2195_c7_45c6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2195_c7_45c6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2195_c7_45c6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2195_c7_45c6]
signal result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2195_c7_45c6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2195_c7_45c6]
signal t8_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2195_c7_45c6]
signal n8_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2198_c11_9acc]
signal BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2198_c7_ea93]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2198_c7_ea93]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2198_c7_ea93]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2198_c7_ea93]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2198_c7_ea93]
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2198_c7_ea93]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2198_c7_ea93]
signal t8_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2198_c7_ea93]
signal n8_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2202_c11_0522]
signal BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2202_c7_8a1c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2202_c7_8a1c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2202_c7_8a1c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2202_c7_8a1c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2202_c7_8a1c]
signal result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2202_c7_8a1c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2202_c7_8a1c]
signal n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2205_c11_26f8]
signal BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2205_c7_37b1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2205_c7_37b1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2205_c7_37b1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2205_c7_37b1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2205_c7_37b1]
signal result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2205_c7_37b1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2205_c7_37b1]
signal n8_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2208_c30_1954]
signal sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2211_c21_d427]
signal BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_return_output : unsigned(0 downto 0);

-- BIN_OP_DIV[uxn_opcodes_h_l2211_c35_7383]
signal BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_left : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_right : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l2211_c21_9c49]
signal MUX_uxn_opcodes_h_l2211_c21_9c49_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2211_c21_9c49_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2211_c21_9c49_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2211_c21_9c49_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2213_c11_1617]
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2213_c7_d361]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2213_c7_d361]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2213_c7_d361]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_641b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77
BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_left,
BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_right,
BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed
result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed
result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_cond,
result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output);

-- t8_MUX_uxn_opcodes_h_l2190_c2_91ed
t8_MUX_uxn_opcodes_h_l2190_c2_91ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2190_c2_91ed_cond,
t8_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue,
t8_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse,
t8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output);

-- n8_MUX_uxn_opcodes_h_l2190_c2_91ed
n8_MUX_uxn_opcodes_h_l2190_c2_91ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2190_c2_91ed_cond,
n8_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue,
n8_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse,
n8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output);

-- printf_uxn_opcodes_h_l2191_c3_4034_uxn_opcodes_h_l2191_c3_4034
printf_uxn_opcodes_h_l2191_c3_4034_uxn_opcodes_h_l2191_c3_4034 : entity work.printf_uxn_opcodes_h_l2191_c3_4034_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2191_c3_4034_uxn_opcodes_h_l2191_c3_4034_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5
BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_left,
BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_right,
BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6
result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6
result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6
result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6
result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output);

-- t8_MUX_uxn_opcodes_h_l2195_c7_45c6
t8_MUX_uxn_opcodes_h_l2195_c7_45c6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2195_c7_45c6_cond,
t8_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue,
t8_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse,
t8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output);

-- n8_MUX_uxn_opcodes_h_l2195_c7_45c6
n8_MUX_uxn_opcodes_h_l2195_c7_45c6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2195_c7_45c6_cond,
n8_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue,
n8_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse,
n8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_left,
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_right,
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93
result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93
result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_cond,
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output);

-- t8_MUX_uxn_opcodes_h_l2198_c7_ea93
t8_MUX_uxn_opcodes_h_l2198_c7_ea93 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2198_c7_ea93_cond,
t8_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue,
t8_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse,
t8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output);

-- n8_MUX_uxn_opcodes_h_l2198_c7_ea93
n8_MUX_uxn_opcodes_h_l2198_c7_ea93 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2198_c7_ea93_cond,
n8_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue,
n8_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse,
n8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522
BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_left,
BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_right,
BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c
result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c
result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c
result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c
result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output);

-- n8_MUX_uxn_opcodes_h_l2202_c7_8a1c
n8_MUX_uxn_opcodes_h_l2202_c7_8a1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond,
n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue,
n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse,
n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8
BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_left,
BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_right,
BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1
result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1
result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1
result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1
result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_cond,
result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1
result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output);

-- n8_MUX_uxn_opcodes_h_l2205_c7_37b1
n8_MUX_uxn_opcodes_h_l2205_c7_37b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2205_c7_37b1_cond,
n8_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue,
n8_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse,
n8_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2208_c30_1954
sp_relative_shift_uxn_opcodes_h_l2208_c30_1954 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_ins,
sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_x,
sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_y,
sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427
BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_left,
BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_right,
BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_return_output);

-- BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383
BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383 : entity work.BIN_OP_DIV_uint8_t_uint8_t_0CLK_a148083c port map (
BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_left,
BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_right,
BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_return_output);

-- MUX_uxn_opcodes_h_l2211_c21_9c49
MUX_uxn_opcodes_h_l2211_c21_9c49 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2211_c21_9c49_cond,
MUX_uxn_opcodes_h_l2211_c21_9c49_iftrue,
MUX_uxn_opcodes_h_l2211_c21_9c49_iffalse,
MUX_uxn_opcodes_h_l2211_c21_9c49_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617
BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_left,
BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_right,
BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361
result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output,
 t8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output,
 n8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output,
 t8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output,
 n8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output,
 t8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output,
 n8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output,
 n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output,
 n8_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output,
 sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_return_output,
 BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_return_output,
 MUX_uxn_opcodes_h_l2211_c21_9c49_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2192_c3_d98b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2190_c2_91ed_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2191_c3_4034_uxn_opcodes_h_l2191_c3_4034_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2196_c3_8410 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2195_c7_45c6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_3587 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2198_c7_ea93_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2203_c3_6874 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2210_c3_3f8e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2205_c7_37b1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2205_c7_37b1_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2211_c21_9c49_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2211_c21_9c49_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2211_c21_9c49_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2211_c21_9c49_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_409b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_1938_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_2712_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_6627_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2213_DUPLICATE_ecdc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2186_l2219_DUPLICATE_77a3_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_3587 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_3587;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2210_c3_3f8e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2210_c3_3f8e;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l2211_c21_9c49_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_y := resize(to_signed(-1, 2), 4);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2192_c3_d98b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2192_c3_d98b;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2196_c3_8410 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2196_c3_8410;
     VAR_sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2203_c3_6874 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2203_c3_6874;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_right := to_unsigned(5, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_left := VAR_phase;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_right := t8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2202_c11_0522] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_left;
     BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_return_output := BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2190_c6_bf77] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_left;
     BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output := BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_1938 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_1938_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2198_c11_9acc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_left;
     BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output := BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2205_c11_26f8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_6627 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_6627_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2213_c11_1617] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_left;
     BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_return_output := BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_return_output;

     -- BIN_OP_DIV[uxn_opcodes_h_l2211_c35_7383] LATENCY=0
     -- Inputs
     BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_left <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_left;
     BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_right <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_right;
     -- Outputs
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_return_output := BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2211_c21_d427] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_left;
     BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_return_output := BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2213_DUPLICATE_ecdc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2213_DUPLICATE_ecdc_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2195_c11_15a5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2208_c30_1954] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_ins;
     sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_x;
     sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_return_output := sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_409b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_409b_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_2712 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_2712_return_output := result.u8_value;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2205_c7_37b1] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2205_c7_37b1_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_MUX_uxn_opcodes_h_l2211_c21_9c49_iffalse := VAR_BIN_OP_DIV_uxn_opcodes_h_l2211_c35_7383_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2190_c2_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2190_c2_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c6_bf77_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2195_c7_45c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2195_c7_45c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2195_c11_15a5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2198_c7_ea93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2198_c7_ea93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_9acc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2202_c11_0522_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2205_c7_37b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2205_c11_26f8_return_output;
     VAR_MUX_uxn_opcodes_h_l2211_c21_9c49_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2211_c21_d427_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_1617_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_6627_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_6627_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_6627_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_6627_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_6627_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2213_DUPLICATE_ecdc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2213_DUPLICATE_ecdc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2213_DUPLICATE_ecdc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2213_DUPLICATE_ecdc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2213_DUPLICATE_ecdc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_409b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_409b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_409b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_409b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_409b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_1938_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_1938_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_1938_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_1938_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2202_l2198_l2195_l2190_l2213_DUPLICATE_1938_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_2712_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_2712_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_2712_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_2712_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2205_l2202_l2198_l2195_l2190_DUPLICATE_2712_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2205_c7_37b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2208_c30_1954_return_output;
     -- MUX[uxn_opcodes_h_l2211_c21_9c49] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2211_c21_9c49_cond <= VAR_MUX_uxn_opcodes_h_l2211_c21_9c49_cond;
     MUX_uxn_opcodes_h_l2211_c21_9c49_iftrue <= VAR_MUX_uxn_opcodes_h_l2211_c21_9c49_iftrue;
     MUX_uxn_opcodes_h_l2211_c21_9c49_iffalse <= VAR_MUX_uxn_opcodes_h_l2211_c21_9c49_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2211_c21_9c49_return_output := MUX_uxn_opcodes_h_l2211_c21_9c49_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2213_c7_d361] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_return_output;

     -- t8_MUX[uxn_opcodes_h_l2198_c7_ea93] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2198_c7_ea93_cond <= VAR_t8_MUX_uxn_opcodes_h_l2198_c7_ea93_cond;
     t8_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue;
     t8_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output := t8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2205_c7_37b1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2213_c7_d361] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2190_c1_9bdd] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_return_output;

     -- n8_MUX[uxn_opcodes_h_l2205_c7_37b1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2205_c7_37b1_cond <= VAR_n8_MUX_uxn_opcodes_h_l2205_c7_37b1_cond;
     n8_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue;
     n8_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output := n8_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2213_c7_d361] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2205_c7_37b1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue := VAR_MUX_uxn_opcodes_h_l2211_c21_9c49_return_output;
     VAR_printf_uxn_opcodes_h_l2191_c3_4034_uxn_opcodes_h_l2191_c3_4034_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2190_c1_9bdd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_d361_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2213_c7_d361_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_d361_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2205_c7_37b1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;

     -- printf_uxn_opcodes_h_l2191_c3_4034[uxn_opcodes_h_l2191_c3_4034] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2191_c3_4034_uxn_opcodes_h_l2191_c3_4034_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2191_c3_4034_uxn_opcodes_h_l2191_c3_4034_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2202_c7_8a1c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2202_c7_8a1c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2202_c7_8a1c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond;
     n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue;
     n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output := n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2205_c7_37b1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;

     -- t8_MUX[uxn_opcodes_h_l2195_c7_45c6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2195_c7_45c6_cond <= VAR_t8_MUX_uxn_opcodes_h_l2195_c7_45c6_cond;
     t8_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue;
     t8_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output := t8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2205_c7_37b1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output := result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2205_c7_37b1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2205_c7_37b1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2202_c7_8a1c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;

     -- t8_MUX[uxn_opcodes_h_l2190_c2_91ed] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2190_c2_91ed_cond <= VAR_t8_MUX_uxn_opcodes_h_l2190_c2_91ed_cond;
     t8_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue;
     t8_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output := t8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2198_c7_ea93] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2202_c7_8a1c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2202_c7_8a1c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2202_c7_8a1c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2198_c7_ea93] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;

     -- n8_MUX[uxn_opcodes_h_l2198_c7_ea93] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2198_c7_ea93_cond <= VAR_n8_MUX_uxn_opcodes_h_l2198_c7_ea93_cond;
     n8_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue;
     n8_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output := n8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2202_c7_8a1c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2198_c7_ea93] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;

     -- n8_MUX[uxn_opcodes_h_l2195_c7_45c6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2195_c7_45c6_cond <= VAR_n8_MUX_uxn_opcodes_h_l2195_c7_45c6_cond;
     n8_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue;
     n8_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output := n8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2195_c7_45c6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2198_c7_ea93] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2195_c7_45c6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2198_c7_ea93] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2198_c7_ea93] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output := result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_ea93_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c2_91ed] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c2_91ed] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output;

     -- n8_MUX[uxn_opcodes_h_l2190_c2_91ed] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2190_c2_91ed_cond <= VAR_n8_MUX_uxn_opcodes_h_l2190_c2_91ed_cond;
     n8_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue;
     n8_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output := n8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2195_c7_45c6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2195_c7_45c6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2195_c7_45c6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2195_c7_45c6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2195_c7_45c6_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2190_c2_91ed] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output := result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c2_91ed] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c2_91ed] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2190_c2_91ed] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2186_l2219_DUPLICATE_77a3 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2186_l2219_DUPLICATE_77a3_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_641b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c2_91ed_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2186_l2219_DUPLICATE_77a3_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2186_l2219_DUPLICATE_77a3_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
