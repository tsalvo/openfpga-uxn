-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity dup2_0CLK_e4095020 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup2_0CLK_e4095020;
architecture arch of dup2_0CLK_e4095020 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2807_c6_30ec]
signal BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2807_c2_fa21]
signal t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2807_c2_fa21]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2807_c2_fa21]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2807_c2_fa21]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2807_c2_fa21]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2807_c2_fa21]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2807_c2_fa21]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2807_c2_fa21]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2807_c2_fa21]
signal result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2807_c2_fa21]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2807_c2_fa21]
signal t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2820_c11_5665]
signal BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2820_c7_2142]
signal t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2820_c7_2142]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2820_c7_2142]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2820_c7_2142]
signal result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2820_c7_2142]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2820_c7_2142]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2820_c7_2142]
signal t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2823_c11_fcdf]
signal BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2823_c7_1cf2]
signal t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2823_c7_1cf2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2823_c7_1cf2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2823_c7_1cf2]
signal result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2823_c7_1cf2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2823_c7_1cf2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2823_c7_1cf2]
signal t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2825_c30_2e73]
signal sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2830_c11_edcd]
signal BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2830_c7_c44f]
signal t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2830_c7_c44f]
signal result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2830_c7_c44f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2830_c7_c44f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2830_c7_c44f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2836_c11_ab05]
signal BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2836_c7_e850]
signal result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2836_c7_e850]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2836_c7_e850]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2840_c11_cac6]
signal BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2840_c7_9ef6]
signal result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2840_c7_9ef6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2840_c7_9ef6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output : unsigned(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a47b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.u8_value := ref_toks_8;
      base.is_vram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec
BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_left,
BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_right,
BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21
t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_cond,
t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue,
t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse,
t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21
result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21
result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21
result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21
result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21
result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21
result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_cond,
result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21
result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21
t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_cond,
t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue,
t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse,
t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665
BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_left,
BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_right,
BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2820_c7_2142
t16_low_MUX_uxn_opcodes_h_l2820_c7_2142 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_cond,
t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue,
t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse,
t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142
result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142
result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142
result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_cond,
result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142
result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2820_c7_2142
t16_high_MUX_uxn_opcodes_h_l2820_c7_2142 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_cond,
t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue,
t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse,
t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf
BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_left,
BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_right,
BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2
t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond,
t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue,
t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse,
t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2
result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2
t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond,
t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue,
t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse,
t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73
sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_ins,
sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_x,
sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_y,
sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd
BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_left,
BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_right,
BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f
t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_cond,
t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue,
t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse,
t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f
result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f
result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05
BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_left,
BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_right,
BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850
result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_cond,
result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850
result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6
BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_left,
BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_right,
BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6
result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6
result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output,
 t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
 t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_return_output,
 t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_return_output,
 t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_return_output,
 t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output,
 t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output,
 sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_return_output,
 t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2812_c3_286f : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2817_c3_faea : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2821_c3_a5bc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2827_c3_9a93 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2832_c3_d9c3 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2833_c3_bbf1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2837_c3_675d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2841_c3_0129 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2840_c7_9ef6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2840_l2807_l2820_DUPLICATE_40b9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2820_l2840_l2836_l2830_l2823_DUPLICATE_6a0d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2830_l2820_DUPLICATE_d222_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2820_l2823_DUPLICATE_02fd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2846_l2803_DUPLICATE_ebd4_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2817_c3_faea := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2817_c3_faea;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2832_c3_d9c3 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2832_c3_d9c3;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2827_c3_9a93 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2827_c3_9a93;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2833_c3_bbf1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2833_c3_bbf1;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_y := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2812_c3_286f := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2812_c3_286f;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2837_c3_675d := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2837_c3_675d;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2821_c3_a5bc := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2821_c3_a5bc;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2841_c3_0129 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2841_c3_0129;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse := t16_high;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse := t16_low;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2820_l2840_l2836_l2830_l2823_DUPLICATE_6a0d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2820_l2840_l2836_l2830_l2823_DUPLICATE_6a0d_return_output := result.is_opc_done;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2807_c2_fa21_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2820_l2823_DUPLICATE_02fd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2820_l2823_DUPLICATE_02fd_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2840_l2807_l2820_DUPLICATE_40b9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2840_l2807_l2820_DUPLICATE_40b9_return_output := result.u8_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2807_c2_fa21_return_output := result.is_ram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2807_c2_fa21_return_output := result.is_stack_index_flipped;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2807_c2_fa21_return_output := result.is_pc_updated;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2830_l2820_DUPLICATE_d222 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2830_l2820_DUPLICATE_d222_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l2825_c30_2e73] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_ins;
     sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_x;
     sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_return_output := sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2840_c11_cac6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2807_c6_30ec] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_left;
     BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output := BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2823_c11_fcdf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_left;
     BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_return_output := BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2836_c11_ab05] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_left;
     BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_return_output := BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2840_c7_9ef6] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2840_c7_9ef6_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2830_c11_edcd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2820_c11_5665] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_left;
     BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_return_output := BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2807_c6_30ec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2820_c11_5665_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_fcdf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2830_c11_edcd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2836_c11_ab05_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2840_c11_cac6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2830_l2820_DUPLICATE_d222_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2830_l2820_DUPLICATE_d222_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2820_l2840_l2836_l2830_l2823_DUPLICATE_6a0d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2820_l2840_l2836_l2830_l2823_DUPLICATE_6a0d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2820_l2840_l2836_l2830_l2823_DUPLICATE_6a0d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2820_l2840_l2836_l2830_l2823_DUPLICATE_6a0d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2820_l2840_l2836_l2830_l2823_DUPLICATE_6a0d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2820_l2823_DUPLICATE_02fd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2820_l2823_DUPLICATE_02fd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2840_l2807_l2820_DUPLICATE_40b9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2840_l2807_l2820_DUPLICATE_40b9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2840_l2807_l2820_DUPLICATE_40b9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2807_c2_fa21_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2807_c2_fa21_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2807_c2_fa21_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2807_c2_fa21_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2840_c7_9ef6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2825_c30_2e73_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2823_c7_1cf2] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond;
     t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output := t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2840_c7_9ef6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2830_c7_c44f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2840_c7_9ef6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2823_c7_1cf2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2830_c7_c44f] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_cond;
     t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output := t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2840_c7_9ef6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2840_c7_9ef6_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2836_c7_e850] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_return_output := result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2823_c7_1cf2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2823_c7_1cf2] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond;
     t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output := t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2820_c7_2142] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2836_c7_e850] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2820_c7_2142] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_cond;
     t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_return_output := t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2836_c7_e850] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2836_c7_e850_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2836_c7_e850_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2836_c7_e850_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;
     -- t16_low_MUX[uxn_opcodes_h_l2820_c7_2142] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_cond;
     t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_return_output := t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2820_c7_2142] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2830_c7_c44f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_cond;
     t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output := t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2830_c7_c44f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2830_c7_c44f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2830_c7_c44f_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2823_c7_1cf2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_cond;
     t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output := t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2823_c7_1cf2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2823_c7_1cf2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_1cf2_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2820_c7_2142] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_return_output := result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2820_c7_2142] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2820_c7_2142] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2820_c7_2142_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output := result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2807_c2_fa21] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2846_l2803_DUPLICATE_ebd4 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2846_l2803_DUPLICATE_ebd4_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a47b(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2807_c2_fa21_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2846_l2803_DUPLICATE_ebd4_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2846_l2803_DUPLICATE_ebd4_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
