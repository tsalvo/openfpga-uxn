-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 42
entity dup_0CLK_6d5e0476 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_6d5e0476;
architecture arch of dup_0CLK_6d5e0476 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l3033_c6_9fa0]
signal BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l3033_c2_75a8]
signal t8_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l3033_c2_75a8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3033_c2_75a8]
signal result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3033_c2_75a8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3033_c2_75a8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3033_c2_75a8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3033_c2_75a8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3038_c11_8afa]
signal BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l3038_c7_832e]
signal t8_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l3038_c7_832e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3038_c7_832e]
signal result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3038_c7_832e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3038_c7_832e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3038_c7_832e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3038_c7_832e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3041_c11_88ea]
signal BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l3041_c7_7364]
signal t8_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l3041_c7_7364]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3041_c7_7364]
signal result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3041_c7_7364]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3041_c7_7364]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3041_c7_7364]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3041_c7_7364]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l3044_c32_cdc0]
signal BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l3044_c32_f75b]
signal BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l3044_c32_609f]
signal MUX_uxn_opcodes_h_l3044_c32_609f_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l3044_c32_609f_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l3044_c32_609f_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l3044_c32_609f_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3046_c11_0620]
signal BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3046_c7_daea]
signal result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3046_c7_daea]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3046_c7_daea]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3046_c7_daea]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3046_c7_daea]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3052_c11_a3dc]
signal BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3052_c7_4d9c]
signal result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3052_c7_4d9c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3052_c7_4d9c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3052_c7_4d9c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3056_c11_adbc]
signal BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3056_c7_43a9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3056_c7_43a9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_value := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_opc_done := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0
BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_left,
BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_right,
BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_return_output);

-- t8_MUX_uxn_opcodes_h_l3033_c2_75a8
t8_MUX_uxn_opcodes_h_l3033_c2_75a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l3033_c2_75a8_cond,
t8_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue,
t8_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse,
t8_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8
result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8
result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_cond,
result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8
result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8
result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8
result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa
BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_left,
BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_right,
BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_return_output);

-- t8_MUX_uxn_opcodes_h_l3038_c7_832e
t8_MUX_uxn_opcodes_h_l3038_c7_832e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l3038_c7_832e_cond,
t8_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue,
t8_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse,
t8_MUX_uxn_opcodes_h_l3038_c7_832e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e
result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e
result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_cond,
result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e
result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e
result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e
result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea
BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_left,
BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_right,
BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_return_output);

-- t8_MUX_uxn_opcodes_h_l3041_c7_7364
t8_MUX_uxn_opcodes_h_l3041_c7_7364 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l3041_c7_7364_cond,
t8_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue,
t8_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse,
t8_MUX_uxn_opcodes_h_l3041_c7_7364_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364
result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364
result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_cond,
result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364
result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364
result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364
result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0
BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_left,
BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_right,
BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b
BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_left,
BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_right,
BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_return_output);

-- MUX_uxn_opcodes_h_l3044_c32_609f
MUX_uxn_opcodes_h_l3044_c32_609f : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l3044_c32_609f_cond,
MUX_uxn_opcodes_h_l3044_c32_609f_iftrue,
MUX_uxn_opcodes_h_l3044_c32_609f_iffalse,
MUX_uxn_opcodes_h_l3044_c32_609f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620
BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_left,
BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_right,
BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea
result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_cond,
result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea
result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea
result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea
result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc
BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_left,
BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_right,
BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c
result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond,
result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc
BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_left,
BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_right,
BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9
result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9
result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_return_output,
 t8_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_return_output,
 t8_MUX_uxn_opcodes_h_l3038_c7_832e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_return_output,
 t8_MUX_uxn_opcodes_h_l3041_c7_7364_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_return_output,
 BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_return_output,
 BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_return_output,
 MUX_uxn_opcodes_h_l3044_c32_609f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3035_c3_449f : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3039_c3_5c21 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3044_c32_609f_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3044_c32_609f_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3044_c32_609f_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3044_c32_609f_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3049_c3_b5f5 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3053_c3_a220 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3038_l3041_l3033_DUPLICATE_c15b_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3038_l3052_l3041_l3033_DUPLICATE_253b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3038_l3033_l3046_DUPLICATE_143c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3041_l3038_l3033_l3056_l3052_DUPLICATE_d9ed_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3041_l3038_l3056_l3052_l3046_DUPLICATE_27f5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3052_l3041_DUPLICATE_0b9f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l3029_l3061_DUPLICATE_dba9_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3035_c3_449f := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3035_c3_449f;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3053_c3_a220 := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3053_c3_a220;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3049_c3_b5f5 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3049_c3_b5f5;
     VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_right := to_unsigned(128, 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3039_c3_5c21 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3039_c3_5c21;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_right := to_unsigned(4, 3);
     VAR_MUX_uxn_opcodes_h_l3044_c32_609f_iftrue := signed(std_logic_vector(resize(to_unsigned(2, 2), 8)));
     VAR_MUX_uxn_opcodes_h_l3044_c32_609f_iffalse := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue := t8;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3052_l3041_DUPLICATE_0b9f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3052_l3041_DUPLICATE_0b9f_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3041_l3038_l3033_l3056_l3052_DUPLICATE_d9ed LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3041_l3038_l3033_l3056_l3052_DUPLICATE_d9ed_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l3056_c11_adbc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_left;
     BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_return_output := BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3038_l3052_l3041_l3033_DUPLICATE_253b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3038_l3052_l3041_l3033_DUPLICATE_253b_return_output := result.stack_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l3046_c11_0620] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_left;
     BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_return_output := BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l3033_c6_9fa0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_left;
     BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_return_output := BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3041_l3038_l3056_l3052_l3046_DUPLICATE_27f5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3041_l3038_l3056_l3052_l3046_DUPLICATE_27f5_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l3041_c11_88ea] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_left;
     BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_return_output := BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3038_l3041_l3033_DUPLICATE_c15b LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3038_l3041_l3033_DUPLICATE_c15b_return_output := result.sp_relative_shift;

     -- BIN_OP_AND[uxn_opcodes_h_l3044_c32_cdc0] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_left;
     BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_return_output := BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l3052_c11_a3dc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_left;
     BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_return_output := BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3038_l3033_l3046_DUPLICATE_143c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3038_l3033_l3046_DUPLICATE_143c_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l3038_c11_8afa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_left;
     BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_return_output := BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_left := VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_cdc0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_9fa0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3038_c7_832e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_8afa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3041_c7_7364_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_88ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_0620_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_a3dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_adbc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3038_l3041_l3033_DUPLICATE_c15b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3038_l3041_l3033_DUPLICATE_c15b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3038_l3041_l3033_DUPLICATE_c15b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3041_l3038_l3056_l3052_l3046_DUPLICATE_27f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3041_l3038_l3056_l3052_l3046_DUPLICATE_27f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3041_l3038_l3056_l3052_l3046_DUPLICATE_27f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3041_l3038_l3056_l3052_l3046_DUPLICATE_27f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3041_l3038_l3056_l3052_l3046_DUPLICATE_27f5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3038_l3033_l3046_DUPLICATE_143c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3038_l3033_l3046_DUPLICATE_143c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3038_l3033_l3046_DUPLICATE_143c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3041_l3038_l3033_l3056_l3052_DUPLICATE_d9ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3041_l3038_l3033_l3056_l3052_DUPLICATE_d9ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3041_l3038_l3033_l3056_l3052_DUPLICATE_d9ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3041_l3038_l3033_l3056_l3052_DUPLICATE_d9ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3041_l3038_l3033_l3056_l3052_DUPLICATE_d9ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3052_l3041_DUPLICATE_0b9f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3052_l3041_DUPLICATE_0b9f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3038_l3052_l3041_l3033_DUPLICATE_253b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3038_l3052_l3041_l3033_DUPLICATE_253b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3038_l3052_l3041_l3033_DUPLICATE_253b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3038_l3052_l3041_l3033_DUPLICATE_253b_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3046_c7_daea] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3056_c7_43a9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l3044_c32_f75b] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_left;
     BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_return_output := BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3056_c7_43a9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3052_c7_4d9c] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output := result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3052_c7_4d9c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output;

     -- t8_MUX[uxn_opcodes_h_l3041_c7_7364] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l3041_c7_7364_cond <= VAR_t8_MUX_uxn_opcodes_h_l3041_c7_7364_cond;
     t8_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue;
     t8_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l3041_c7_7364_return_output := t8_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l3044_c32_609f_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_f75b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_daea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_43a9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3041_c7_7364] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;

     -- t8_MUX[uxn_opcodes_h_l3038_c7_832e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l3038_c7_832e_cond <= VAR_t8_MUX_uxn_opcodes_h_l3038_c7_832e_cond;
     t8_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue;
     t8_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l3038_c7_832e_return_output := t8_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3052_c7_4d9c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3046_c7_daea] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_return_output := result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3046_c7_daea] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_return_output;

     -- MUX[uxn_opcodes_h_l3044_c32_609f] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l3044_c32_609f_cond <= VAR_MUX_uxn_opcodes_h_l3044_c32_609f_cond;
     MUX_uxn_opcodes_h_l3044_c32_609f_iftrue <= VAR_MUX_uxn_opcodes_h_l3044_c32_609f_iftrue;
     MUX_uxn_opcodes_h_l3044_c32_609f_iffalse <= VAR_MUX_uxn_opcodes_h_l3044_c32_609f_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l3044_c32_609f_return_output := MUX_uxn_opcodes_h_l3044_c32_609f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3052_c7_4d9c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue := VAR_MUX_uxn_opcodes_h_l3044_c32_609f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_4d9c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_daea_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_daea_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;
     -- t8_MUX[uxn_opcodes_h_l3033_c2_75a8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l3033_c2_75a8_cond <= VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75a8_cond;
     t8_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue;
     t8_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output := t8_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l3041_c7_7364] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3041_c7_7364] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_return_output := result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3038_c7_832e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3041_c7_7364] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3046_c7_daea] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3046_c7_daea] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_daea_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_daea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3038_c7_832e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3041_c7_7364] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l3038_c7_832e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3033_c2_75a8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3041_c7_7364] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3038_c7_832e] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_return_output := result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_7364_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l3038_c7_832e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l3033_c2_75a8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3033_c2_75a8] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output := result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3038_c7_832e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3033_c2_75a8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_832e_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l3033_c2_75a8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3033_c2_75a8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l3029_l3061_DUPLICATE_dba9 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l3029_l3061_DUPLICATE_dba9_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75a8_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l3029_l3061_DUPLICATE_dba9_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l3029_l3061_DUPLICATE_dba9_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
