-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity ovr_0CLK_61914e8d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ovr_0CLK_61914e8d;
architecture arch of ovr_0CLK_61914e8d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l297_c6_9382]
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l297_c2_aae7]
signal n8_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l297_c2_aae7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l297_c2_aae7]
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l297_c2_aae7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l297_c2_aae7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l297_c2_aae7]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l297_c2_aae7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l297_c2_aae7]
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l297_c2_aae7]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l297_c2_aae7]
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l297_c2_aae7]
signal t8_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l310_c11_3205]
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l310_c7_7f93]
signal n8_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l310_c7_7f93]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l310_c7_7f93]
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l310_c7_7f93]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l310_c7_7f93]
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l310_c7_7f93]
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l310_c7_7f93]
signal t8_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l313_c11_9d18]
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l313_c7_5d33]
signal n8_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l313_c7_5d33]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l313_c7_5d33]
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l313_c7_5d33]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l313_c7_5d33]
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l313_c7_5d33]
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l313_c7_5d33]
signal t8_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l315_c30_63ca]
signal sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l320_c11_572f]
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l320_c7_c507]
signal n8_MUX_uxn_opcodes_h_l320_c7_c507_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_c507_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_c507_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_c507_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l320_c7_c507]
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l320_c7_c507]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l320_c7_c507]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l320_c7_c507]
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l326_c11_5437]
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l326_c7_d4dc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l326_c7_d4dc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l326_c7_d4dc]
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_04b4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382
BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_left,
BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_right,
BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output);

-- n8_MUX_uxn_opcodes_h_l297_c2_aae7
n8_MUX_uxn_opcodes_h_l297_c2_aae7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l297_c2_aae7_cond,
n8_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue,
n8_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse,
n8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7
result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_cond,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_return_output);

-- t8_MUX_uxn_opcodes_h_l297_c2_aae7
t8_MUX_uxn_opcodes_h_l297_c2_aae7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l297_c2_aae7_cond,
t8_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue,
t8_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse,
t8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205
BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_left,
BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_right,
BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_return_output);

-- n8_MUX_uxn_opcodes_h_l310_c7_7f93
n8_MUX_uxn_opcodes_h_l310_c7_7f93 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l310_c7_7f93_cond,
n8_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue,
n8_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse,
n8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93
result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_cond,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_return_output);

-- t8_MUX_uxn_opcodes_h_l310_c7_7f93
t8_MUX_uxn_opcodes_h_l310_c7_7f93 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l310_c7_7f93_cond,
t8_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue,
t8_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse,
t8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18
BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_left,
BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_right,
BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_return_output);

-- n8_MUX_uxn_opcodes_h_l313_c7_5d33
n8_MUX_uxn_opcodes_h_l313_c7_5d33 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l313_c7_5d33_cond,
n8_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue,
n8_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse,
n8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33
result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_cond,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_return_output);

-- t8_MUX_uxn_opcodes_h_l313_c7_5d33
t8_MUX_uxn_opcodes_h_l313_c7_5d33 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l313_c7_5d33_cond,
t8_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue,
t8_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse,
t8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output);

-- sp_relative_shift_uxn_opcodes_h_l315_c30_63ca
sp_relative_shift_uxn_opcodes_h_l315_c30_63ca : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_ins,
sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_x,
sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_y,
sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f
BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_left,
BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_right,
BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_return_output);

-- n8_MUX_uxn_opcodes_h_l320_c7_c507
n8_MUX_uxn_opcodes_h_l320_c7_c507 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l320_c7_c507_cond,
n8_MUX_uxn_opcodes_h_l320_c7_c507_iftrue,
n8_MUX_uxn_opcodes_h_l320_c7_c507_iffalse,
n8_MUX_uxn_opcodes_h_l320_c7_c507_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507
result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_cond,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437
BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_left,
BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_right,
BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc
result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_cond,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output,
 n8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
 t8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_return_output,
 n8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_return_output,
 t8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_return_output,
 n8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_return_output,
 t8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output,
 sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_return_output,
 n8_MUX_uxn_opcodes_h_l320_c7_c507_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_247b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_d21c : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_aae7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_4005 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_7f93_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_c507_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_484a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_5d33_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_c507_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_c507_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_c507_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l322_c3_addb : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_1eeb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_6a9e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_d4dc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l310_l326_l297_DUPLICATE_c88d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l310_l320_DUPLICATE_9bae_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_8de5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_802d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l332_l293_DUPLICATE_5bfb_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_4005 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_4005;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_right := to_unsigned(2, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_d21c := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_d21c;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_1eeb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_1eeb;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_247b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_247b;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l322_c3_addb := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l322_c3_addb;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_484a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_484a;
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_6a9e := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_6a9e;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_right := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_right := to_unsigned(4, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_c507_iffalse := n8;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_c507_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse := t8;
     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_aae7_return_output := result.is_stack_index_flipped;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l326_c7_d4dc] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_d4dc_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l313_c11_9d18] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_left;
     BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_return_output := BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_aae7_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l326_c11_5437] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_left;
     BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_return_output := BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_aae7_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l297_c6_9382] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_left;
     BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output := BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_aae7_return_output := result.is_vram_write;

     -- sp_relative_shift[uxn_opcodes_h_l315_c30_63ca] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_ins;
     sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_x <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_x;
     sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_y <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_return_output := sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_802d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_802d_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_8de5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_8de5_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l320_c11_572f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_left;
     BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_return_output := BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l310_l320_DUPLICATE_9bae LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l310_l320_DUPLICATE_9bae_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l310_l326_l297_DUPLICATE_c88d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l310_l326_l297_DUPLICATE_c88d_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l310_c11_3205] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_left;
     BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_return_output := BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_aae7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_aae7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_9382_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_7f93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_7f93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_3205_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_5d33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_5d33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_9d18_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_c507_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_572f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5437_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l310_l320_DUPLICATE_9bae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l310_l320_DUPLICATE_9bae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_8de5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_8de5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_8de5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_8de5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_802d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_802d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l310_l326_l297_DUPLICATE_c88d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l310_l326_l297_DUPLICATE_c88d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l310_l326_l297_DUPLICATE_c88d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_aae7_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_aae7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_aae7_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_aae7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_d4dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_63ca_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l326_c7_d4dc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output := result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l313_c7_5d33] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l326_c7_d4dc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output;

     -- n8_MUX[uxn_opcodes_h_l320_c7_c507] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l320_c7_c507_cond <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_c507_cond;
     n8_MUX_uxn_opcodes_h_l320_c7_c507_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_c507_iftrue;
     n8_MUX_uxn_opcodes_h_l320_c7_c507_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_c507_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_c507_return_output := n8_MUX_uxn_opcodes_h_l320_c7_c507_return_output;

     -- t8_MUX[uxn_opcodes_h_l313_c7_5d33] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l313_c7_5d33_cond <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_5d33_cond;
     t8_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue;
     t8_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output := t8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l320_c7_c507] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l326_c7_d4dc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse := VAR_n8_MUX_uxn_opcodes_h_l320_c7_c507_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_c507_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_d4dc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse := VAR_t8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l320_c7_c507] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_cond;
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_return_output := result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l310_c7_7f93] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l320_c7_c507] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_return_output;

     -- t8_MUX[uxn_opcodes_h_l310_c7_7f93] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l310_c7_7f93_cond <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_7f93_cond;
     t8_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue;
     t8_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output := t8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;

     -- n8_MUX[uxn_opcodes_h_l313_c7_5d33] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l313_c7_5d33_cond <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_5d33_cond;
     n8_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue;
     n8_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output := n8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l320_c7_c507] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l313_c7_5d33] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse := VAR_n8_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_c507_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_c507_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_c507_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse := VAR_t8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;
     -- t8_MUX[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l297_c2_aae7_cond <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_aae7_cond;
     t8_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue;
     t8_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output := t8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l313_c7_5d33] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_cond;
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_return_output := result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l310_c7_7f93] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;

     -- n8_MUX[uxn_opcodes_h_l310_c7_7f93] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l310_c7_7f93_cond <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_7f93_cond;
     n8_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue;
     n8_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output := n8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l313_c7_5d33] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l313_c7_5d33] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse := VAR_n8_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_5d33_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output;
     -- n8_MUX[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l297_c2_aae7_cond <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_aae7_cond;
     n8_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue;
     n8_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output := n8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l310_c7_7f93] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l310_c7_7f93] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l310_c7_7f93] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_cond;
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_return_output := result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l297_c2_aae7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_7f93_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_return_output := result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l297_c2_aae7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l332_l293_DUPLICATE_5bfb LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l332_l293_DUPLICATE_5bfb_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_04b4(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_aae7_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_aae7_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l332_l293_DUPLICATE_5bfb_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l332_l293_DUPLICATE_5bfb_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
