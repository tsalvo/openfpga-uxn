-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity eor_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor_0CLK_f62d646e;
architecture arch of eor_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1138_c6_ca11]
signal BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1138_c1_318e]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1138_c2_eb95]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1138_c2_eb95]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1138_c2_eb95]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1138_c2_eb95]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1138_c2_eb95]
signal result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1138_c2_eb95]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1138_c2_eb95]
signal t8_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1138_c2_eb95]
signal n8_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1139_c3_8dd1[uxn_opcodes_h_l1139_c3_8dd1]
signal printf_uxn_opcodes_h_l1139_c3_8dd1_uxn_opcodes_h_l1139_c3_8dd1_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1143_c11_6cf6]
signal BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1143_c7_6f60]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1143_c7_6f60]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1143_c7_6f60]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1143_c7_6f60]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1143_c7_6f60]
signal result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1143_c7_6f60]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1143_c7_6f60]
signal t8_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1143_c7_6f60]
signal n8_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1146_c11_8575]
signal BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1146_c7_6819]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1146_c7_6819]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1146_c7_6819]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1146_c7_6819]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1146_c7_6819]
signal result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1146_c7_6819]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1146_c7_6819]
signal t8_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1146_c7_6819]
signal n8_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1150_c11_d4a5]
signal BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1150_c7_9067]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1150_c7_9067]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1150_c7_9067]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1150_c7_9067]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1150_c7_9067]
signal result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1150_c7_9067]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1150_c7_9067]
signal n8_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1153_c11_c559]
signal BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1153_c7_ecd2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1153_c7_ecd2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1153_c7_ecd2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1153_c7_ecd2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1153_c7_ecd2]
signal result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1153_c7_ecd2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1153_c7_ecd2]
signal n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1156_c30_7269]
signal sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_return_output : signed(3 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1159_c21_d325]
signal BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_left : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_right : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1161_c11_3069]
signal BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1161_c7_45b9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1161_c7_45b9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1161_c7_45b9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_641b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11
BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_left,
BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_right,
BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95
result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95
result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95
result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95
result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_cond,
result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95
result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output);

-- t8_MUX_uxn_opcodes_h_l1138_c2_eb95
t8_MUX_uxn_opcodes_h_l1138_c2_eb95 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1138_c2_eb95_cond,
t8_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue,
t8_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse,
t8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output);

-- n8_MUX_uxn_opcodes_h_l1138_c2_eb95
n8_MUX_uxn_opcodes_h_l1138_c2_eb95 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1138_c2_eb95_cond,
n8_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue,
n8_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse,
n8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output);

-- printf_uxn_opcodes_h_l1139_c3_8dd1_uxn_opcodes_h_l1139_c3_8dd1
printf_uxn_opcodes_h_l1139_c3_8dd1_uxn_opcodes_h_l1139_c3_8dd1 : entity work.printf_uxn_opcodes_h_l1139_c3_8dd1_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1139_c3_8dd1_uxn_opcodes_h_l1139_c3_8dd1_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6
BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_left,
BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_right,
BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60
result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60
result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60
result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60
result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_cond,
result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60
result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output);

-- t8_MUX_uxn_opcodes_h_l1143_c7_6f60
t8_MUX_uxn_opcodes_h_l1143_c7_6f60 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1143_c7_6f60_cond,
t8_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue,
t8_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse,
t8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output);

-- n8_MUX_uxn_opcodes_h_l1143_c7_6f60
n8_MUX_uxn_opcodes_h_l1143_c7_6f60 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1143_c7_6f60_cond,
n8_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue,
n8_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse,
n8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575
BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_left,
BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_right,
BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819
result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819
result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819
result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819
result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_cond,
result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819
result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output);

-- t8_MUX_uxn_opcodes_h_l1146_c7_6819
t8_MUX_uxn_opcodes_h_l1146_c7_6819 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1146_c7_6819_cond,
t8_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue,
t8_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse,
t8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output);

-- n8_MUX_uxn_opcodes_h_l1146_c7_6819
n8_MUX_uxn_opcodes_h_l1146_c7_6819 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1146_c7_6819_cond,
n8_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue,
n8_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse,
n8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5
BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_left,
BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_right,
BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067
result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067
result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067
result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067
result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_cond,
result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067
result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output);

-- n8_MUX_uxn_opcodes_h_l1150_c7_9067
n8_MUX_uxn_opcodes_h_l1150_c7_9067 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1150_c7_9067_cond,
n8_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue,
n8_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse,
n8_MUX_uxn_opcodes_h_l1150_c7_9067_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559
BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_left,
BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_right,
BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2
result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2
result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2
result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2
result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output);

-- n8_MUX_uxn_opcodes_h_l1153_c7_ecd2
n8_MUX_uxn_opcodes_h_l1153_c7_ecd2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond,
n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue,
n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse,
n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1156_c30_7269
sp_relative_shift_uxn_opcodes_h_l1156_c30_7269 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_ins,
sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_x,
sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_y,
sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325
BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325 : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_left,
BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_right,
BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069
BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_left,
BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_right,
BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9
result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9
result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9
result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output,
 t8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output,
 n8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output,
 t8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output,
 n8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output,
 t8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output,
 n8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output,
 n8_MUX_uxn_opcodes_h_l1150_c7_9067_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output,
 n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output,
 sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1140_c3_a099 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1138_c2_eb95_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1139_c3_8dd1_uxn_opcodes_h_l1139_c3_8dd1_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1144_c3_b080 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1143_c7_6f60_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1148_c3_34b7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1150_c7_9067_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1146_c7_6819_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1151_c3_b636 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1150_c7_9067_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1158_c3_665c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1153_c7_ecd2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_1141_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_eca7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_fa3f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_cf66_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1143_l1161_l1153_l1150_l1146_DUPLICATE_0456_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1167_l1134_DUPLICATE_d567_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1144_c3_b080 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1144_c3_b080;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1158_c3_665c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1158_c3_665c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1148_c3_34b7 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1148_c3_34b7;
     VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1140_c3_a099 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1140_c3_a099;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_iffalse := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1151_c3_b636 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1151_c3_b636;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_right := to_unsigned(5, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1143_c11_6cf6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_left;
     BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output := BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1150_c11_d4a5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_1141 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_1141_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_fa3f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_fa3f_return_output := result.u8_value;

     -- BIN_OP_XOR[uxn_opcodes_h_l1159_c21_d325] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_left;
     BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_return_output := BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1161_c11_3069] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_left;
     BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_return_output := BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1143_l1161_l1153_l1150_l1146_DUPLICATE_0456 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1143_l1161_l1153_l1150_l1146_DUPLICATE_0456_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_eca7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_eca7_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1146_c11_8575] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_left;
     BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output := BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1156_c30_7269] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_ins;
     sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_x;
     sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_return_output := sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1138_c6_ca11] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_left;
     BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output := BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1153_c11_c559] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_left;
     BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_return_output := BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1153_c7_ecd2] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1153_c7_ecd2_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_cf66 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_cf66_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1138_c2_eb95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1138_c2_eb95_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1138_c6_ca11_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1143_c7_6f60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1143_c7_6f60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1143_c11_6cf6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1146_c7_6819_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1146_c7_6819_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1146_c11_8575_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1150_c7_9067_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_d4a5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_c559_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_3069_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1159_c21_d325_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_cf66_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_cf66_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_cf66_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_cf66_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_cf66_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1143_l1161_l1153_l1150_l1146_DUPLICATE_0456_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1143_l1161_l1153_l1150_l1146_DUPLICATE_0456_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1143_l1161_l1153_l1150_l1146_DUPLICATE_0456_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1143_l1161_l1153_l1150_l1146_DUPLICATE_0456_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1143_l1161_l1153_l1150_l1146_DUPLICATE_0456_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_1141_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_1141_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_1141_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_1141_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_1141_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_eca7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_eca7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_eca7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_eca7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1143_l1138_l1161_l1150_l1146_DUPLICATE_eca7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_fa3f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_fa3f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_fa3f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_fa3f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1143_l1138_l1153_l1150_l1146_DUPLICATE_fa3f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1153_c7_ecd2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_7269_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1161_c7_45b9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output;

     -- t8_MUX[uxn_opcodes_h_l1146_c7_6819] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1146_c7_6819_cond <= VAR_t8_MUX_uxn_opcodes_h_l1146_c7_6819_cond;
     t8_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue;
     t8_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output := t8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;

     -- n8_MUX[uxn_opcodes_h_l1153_c7_ecd2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond <= VAR_n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond;
     n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue;
     n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output := n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1161_c7_45b9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1153_c7_ecd2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1161_c7_45b9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1153_c7_ecd2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1153_c7_ecd2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1138_c1_318e] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l1139_c3_8dd1_uxn_opcodes_h_l1139_c3_8dd1_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1138_c1_318e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_45b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1150_c7_9067] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1153_c7_ecd2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;

     -- t8_MUX[uxn_opcodes_h_l1143_c7_6f60] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1143_c7_6f60_cond <= VAR_t8_MUX_uxn_opcodes_h_l1143_c7_6f60_cond;
     t8_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue;
     t8_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output := t8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1150_c7_9067] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1153_c7_ecd2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;

     -- printf_uxn_opcodes_h_l1139_c3_8dd1[uxn_opcodes_h_l1139_c3_8dd1] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1139_c3_8dd1_uxn_opcodes_h_l1139_c3_8dd1_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1139_c3_8dd1_uxn_opcodes_h_l1139_c3_8dd1_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l1150_c7_9067] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_return_output := result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1153_c7_ecd2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;

     -- n8_MUX[uxn_opcodes_h_l1150_c7_9067] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1150_c7_9067_cond <= VAR_n8_MUX_uxn_opcodes_h_l1150_c7_9067_cond;
     n8_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue;
     n8_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1150_c7_9067_return_output := n8_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_ecd2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;
     -- n8_MUX[uxn_opcodes_h_l1146_c7_6819] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1146_c7_6819_cond <= VAR_n8_MUX_uxn_opcodes_h_l1146_c7_6819_cond;
     n8_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue;
     n8_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output := n8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1146_c7_6819] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1150_c7_9067] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1150_c7_9067] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1146_c7_6819] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;

     -- t8_MUX[uxn_opcodes_h_l1138_c2_eb95] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1138_c2_eb95_cond <= VAR_t8_MUX_uxn_opcodes_h_l1138_c2_eb95_cond;
     t8_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue;
     t8_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output := t8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1146_c7_6819] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_return_output := result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1150_c7_9067] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_9067_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output;
     -- n8_MUX[uxn_opcodes_h_l1143_c7_6f60] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1143_c7_6f60_cond <= VAR_n8_MUX_uxn_opcodes_h_l1143_c7_6f60_cond;
     n8_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue;
     n8_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output := n8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1146_c7_6819] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1143_c7_6f60] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1146_c7_6819] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1143_c7_6f60] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1146_c7_6819] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1143_c7_6f60] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output := result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1146_c7_6819_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1138_c2_eb95] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1138_c2_eb95] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output := result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1143_c7_6f60] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;

     -- n8_MUX[uxn_opcodes_h_l1138_c2_eb95] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1138_c2_eb95_cond <= VAR_n8_MUX_uxn_opcodes_h_l1138_c2_eb95_cond;
     n8_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue;
     n8_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output := n8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1138_c2_eb95] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1143_c7_6f60] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1143_c7_6f60] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1143_c7_6f60_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1138_c2_eb95] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1138_c2_eb95] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1138_c2_eb95] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1167_l1134_DUPLICATE_d567 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1167_l1134_DUPLICATE_d567_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_641b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1138_c2_eb95_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1167_l1134_DUPLICATE_d567_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1167_l1134_DUPLICATE_d567_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
