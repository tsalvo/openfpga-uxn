-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 46
entity div_0CLK_a35230ee is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end div_0CLK_a35230ee;
architecture arch of div_0CLK_a35230ee is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1945_c6_9fa5]
signal BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1945_c1_deb7]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1945_c2_912c]
signal n8_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1945_c2_912c]
signal t8_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1945_c2_912c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1945_c2_912c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1945_c2_912c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1945_c2_912c]
signal result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1945_c2_912c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1945_c2_912c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l1946_c3_02e7[uxn_opcodes_h_l1946_c3_02e7]
signal printf_uxn_opcodes_h_l1946_c3_02e7_uxn_opcodes_h_l1946_c3_02e7_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1950_c11_21b3]
signal BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1950_c7_8fe5]
signal n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1950_c7_8fe5]
signal t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1950_c7_8fe5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1950_c7_8fe5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1950_c7_8fe5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1950_c7_8fe5]
signal result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1950_c7_8fe5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1950_c7_8fe5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1953_c11_98ae]
signal BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1953_c7_7099]
signal n8_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1953_c7_7099]
signal t8_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1953_c7_7099]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1953_c7_7099]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1953_c7_7099]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1953_c7_7099]
signal result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1953_c7_7099]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1953_c7_7099]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1956_c11_4451]
signal BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1956_c7_3888]
signal n8_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1956_c7_3888]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1956_c7_3888]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1956_c7_3888]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1956_c7_3888]
signal result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1956_c7_3888]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1956_c7_3888]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1959_c30_62b0]
signal sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1962_c21_4563]
signal BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_return_output : unsigned(0 downto 0);

-- BIN_OP_DIV[uxn_opcodes_h_l1962_c35_2f48]
signal BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_left : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_right : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l1962_c21_f4ec]
signal MUX_uxn_opcodes_h_l1962_c21_f4ec_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1962_c21_f4ec_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1962_c21_f4ec_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1962_c21_f4ec_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1964_c11_2f0e]
signal BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1964_c7_7b44]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1964_c7_7b44]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1964_c7_7b44]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c551( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5
BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_left,
BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_right,
BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_return_output);

-- n8_MUX_uxn_opcodes_h_l1945_c2_912c
n8_MUX_uxn_opcodes_h_l1945_c2_912c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1945_c2_912c_cond,
n8_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue,
n8_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse,
n8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output);

-- t8_MUX_uxn_opcodes_h_l1945_c2_912c
t8_MUX_uxn_opcodes_h_l1945_c2_912c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1945_c2_912c_cond,
t8_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue,
t8_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse,
t8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c
result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c
result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c
result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c
result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output);

-- printf_uxn_opcodes_h_l1946_c3_02e7_uxn_opcodes_h_l1946_c3_02e7
printf_uxn_opcodes_h_l1946_c3_02e7_uxn_opcodes_h_l1946_c3_02e7 : entity work.printf_uxn_opcodes_h_l1946_c3_02e7_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1946_c3_02e7_uxn_opcodes_h_l1946_c3_02e7_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3
BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_left,
BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_right,
BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output);

-- n8_MUX_uxn_opcodes_h_l1950_c7_8fe5
n8_MUX_uxn_opcodes_h_l1950_c7_8fe5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond,
n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue,
n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse,
n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output);

-- t8_MUX_uxn_opcodes_h_l1950_c7_8fe5
t8_MUX_uxn_opcodes_h_l1950_c7_8fe5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond,
t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue,
t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse,
t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5
result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5
result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5
result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5
result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae
BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_left,
BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_right,
BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output);

-- n8_MUX_uxn_opcodes_h_l1953_c7_7099
n8_MUX_uxn_opcodes_h_l1953_c7_7099 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1953_c7_7099_cond,
n8_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue,
n8_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse,
n8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output);

-- t8_MUX_uxn_opcodes_h_l1953_c7_7099
t8_MUX_uxn_opcodes_h_l1953_c7_7099 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1953_c7_7099_cond,
t8_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue,
t8_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse,
t8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099
result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_cond,
result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099
result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451
BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_left,
BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_right,
BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_return_output);

-- n8_MUX_uxn_opcodes_h_l1956_c7_3888
n8_MUX_uxn_opcodes_h_l1956_c7_3888 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1956_c7_3888_cond,
n8_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue,
n8_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse,
n8_MUX_uxn_opcodes_h_l1956_c7_3888_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888
result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888
result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888
result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_cond,
result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888
result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888
result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0
sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_ins,
sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_x,
sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_y,
sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563
BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_left,
BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_right,
BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_return_output);

-- BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48
BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48 : entity work.BIN_OP_DIV_uint8_t_uint8_t_0CLK_a148083c port map (
BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_left,
BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_right,
BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_return_output);

-- MUX_uxn_opcodes_h_l1962_c21_f4ec
MUX_uxn_opcodes_h_l1962_c21_f4ec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1962_c21_f4ec_cond,
MUX_uxn_opcodes_h_l1962_c21_f4ec_iftrue,
MUX_uxn_opcodes_h_l1962_c21_f4ec_iffalse,
MUX_uxn_opcodes_h_l1962_c21_f4ec_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e
BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_left,
BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_right,
BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_return_output,
 n8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output,
 t8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output,
 n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output,
 t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output,
 n8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output,
 t8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_return_output,
 n8_MUX_uxn_opcodes_h_l1956_c7_3888_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output,
 sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_return_output,
 BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_return_output,
 MUX_uxn_opcodes_h_l1962_c21_f4ec_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1947_c3_a133 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1946_c3_02e7_uxn_opcodes_h_l1946_c3_02e7_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1951_c3_043e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1961_c3_dc91 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1962_c21_f4ec_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1962_c21_f4ec_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1962_c21_f4ec_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1962_c21_f4ec_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_e280_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_6e99_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_f6e1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_6e07_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1953_l1956_l1950_l1964_DUPLICATE_84bb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1953_l1956_DUPLICATE_64c2_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l1970_l1941_DUPLICATE_c5f1_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_iffalse := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1962_c21_f4ec_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1961_c3_dc91 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1961_c3_dc91;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1947_c3_a133 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1947_c3_a133;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1951_c3_043e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1951_c3_043e;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_left := VAR_phase;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_right := t8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_f6e1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_f6e1_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1945_c6_9fa5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1962_c21_4563] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_left;
     BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_return_output := BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1953_l1956_l1950_l1964_DUPLICATE_84bb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1953_l1956_l1950_l1964_DUPLICATE_84bb_return_output := result.is_opc_done;

     -- BIN_OP_DIV[uxn_opcodes_h_l1962_c35_2f48] LATENCY=0
     -- Inputs
     BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_left <= VAR_BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_left;
     BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_right <= VAR_BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_right;
     -- Outputs
     VAR_BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_return_output := BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1959_c30_62b0] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_ins;
     sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_x;
     sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_return_output := sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_6e99 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_6e99_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1956_c11_4451] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_left;
     BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_return_output := BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1950_c11_21b3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1953_c11_98ae] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_left;
     BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output := BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1964_c11_2f0e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_6e07 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_6e07_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_e280 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_e280_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1953_l1956_DUPLICATE_64c2 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1953_l1956_DUPLICATE_64c2_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_MUX_uxn_opcodes_h_l1962_c21_f4ec_iffalse := VAR_BIN_OP_DIV_uxn_opcodes_h_l1962_c35_2f48_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1945_c2_912c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1945_c2_912c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1945_c6_9fa5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1950_c11_21b3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1953_c7_7099_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1953_c7_7099_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c11_98ae_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1956_c7_3888_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1956_c11_4451_return_output;
     VAR_MUX_uxn_opcodes_h_l1962_c21_f4ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1962_c21_4563_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_2f0e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_6e99_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_6e99_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_6e99_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_6e99_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1953_l1956_l1950_l1964_DUPLICATE_84bb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1953_l1956_l1950_l1964_DUPLICATE_84bb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1953_l1956_l1950_l1964_DUPLICATE_84bb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1953_l1956_l1950_l1964_DUPLICATE_84bb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_6e07_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_6e07_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_6e07_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_6e07_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_e280_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_e280_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_e280_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1953_l1945_l1950_l1964_DUPLICATE_e280_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1953_l1956_DUPLICATE_64c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1953_l1956_DUPLICATE_64c2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_f6e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_f6e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_f6e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1953_l1945_l1956_l1950_DUPLICATE_f6e1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1959_c30_62b0_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1945_c1_deb7] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_return_output;

     -- n8_MUX[uxn_opcodes_h_l1956_c7_3888] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1956_c7_3888_cond <= VAR_n8_MUX_uxn_opcodes_h_l1956_c7_3888_cond;
     n8_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue;
     n8_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1956_c7_3888_return_output := n8_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1964_c7_7b44] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1956_c7_3888] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1956_c7_3888] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;

     -- MUX[uxn_opcodes_h_l1962_c21_f4ec] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1962_c21_f4ec_cond <= VAR_MUX_uxn_opcodes_h_l1962_c21_f4ec_cond;
     MUX_uxn_opcodes_h_l1962_c21_f4ec_iftrue <= VAR_MUX_uxn_opcodes_h_l1962_c21_f4ec_iftrue;
     MUX_uxn_opcodes_h_l1962_c21_f4ec_iffalse <= VAR_MUX_uxn_opcodes_h_l1962_c21_f4ec_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1962_c21_f4ec_return_output := MUX_uxn_opcodes_h_l1962_c21_f4ec_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1964_c7_7b44] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output;

     -- t8_MUX[uxn_opcodes_h_l1953_c7_7099] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1953_c7_7099_cond <= VAR_t8_MUX_uxn_opcodes_h_l1953_c7_7099_cond;
     t8_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue;
     t8_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output := t8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1964_c7_7b44] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue := VAR_MUX_uxn_opcodes_h_l1962_c21_f4ec_return_output;
     VAR_printf_uxn_opcodes_h_l1946_c3_02e7_uxn_opcodes_h_l1946_c3_02e7_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1945_c1_deb7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_7b44_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1953_c7_7099] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1956_c7_3888] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_return_output := result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1953_c7_7099] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;

     -- t8_MUX[uxn_opcodes_h_l1950_c7_8fe5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond <= VAR_t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond;
     t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue;
     t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output := t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1956_c7_3888] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;

     -- printf_uxn_opcodes_h_l1946_c3_02e7[uxn_opcodes_h_l1946_c3_02e7] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1946_c3_02e7_uxn_opcodes_h_l1946_c3_02e7_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1946_c3_02e7_uxn_opcodes_h_l1946_c3_02e7_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1956_c7_3888] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;

     -- n8_MUX[uxn_opcodes_h_l1953_c7_7099] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1953_c7_7099_cond <= VAR_n8_MUX_uxn_opcodes_h_l1953_c7_7099_cond;
     n8_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue;
     n8_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output := n8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1956_c7_3888] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1956_c7_3888_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1953_c7_7099] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;

     -- t8_MUX[uxn_opcodes_h_l1945_c2_912c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1945_c2_912c_cond <= VAR_t8_MUX_uxn_opcodes_h_l1945_c2_912c_cond;
     t8_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue;
     t8_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output := t8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1953_c7_7099] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1953_c7_7099] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;

     -- n8_MUX[uxn_opcodes_h_l1950_c7_8fe5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond <= VAR_n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond;
     n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue;
     n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output := n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1953_c7_7099] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_return_output := result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1950_c7_8fe5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1950_c7_8fe5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c7_7099_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1945_c2_912c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1945_c2_912c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1950_c7_8fe5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1950_c7_8fe5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;

     -- n8_MUX[uxn_opcodes_h_l1945_c2_912c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1945_c2_912c_cond <= VAR_n8_MUX_uxn_opcodes_h_l1945_c2_912c_cond;
     n8_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue;
     n8_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output := n8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1950_c7_8fe5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1950_c7_8fe5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1945_c2_912c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1950_c7_8fe5_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1945_c2_912c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1945_c2_912c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1945_c2_912c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1945_c2_912c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l1970_l1941_DUPLICATE_c5f1 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l1970_l1941_DUPLICATE_c5f1_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c551(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1945_c2_912c_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1945_c2_912c_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1945_c2_912c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1945_c2_912c_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1945_c2_912c_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l1970_l1941_DUPLICATE_c5f1_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l1970_l1941_DUPLICATE_c5f1_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
