-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 46
entity ovr_0CLK_9159c4aa is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ovr_0CLK_9159c4aa;
architecture arch of ovr_0CLK_9159c4aa is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l286_c6_85cf]
signal BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l286_c1_1890]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l286_c2_7f12]
signal n8_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l286_c2_7f12]
signal t8_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l286_c2_7f12]
signal result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l286_c2_7f12]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l286_c2_7f12]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l286_c2_7f12]
signal result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l286_c2_7f12]
signal result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l286_c2_7f12]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l287_c3_ed90[uxn_opcodes_h_l287_c3_ed90]
signal printf_uxn_opcodes_h_l287_c3_ed90_uxn_opcodes_h_l287_c3_ed90_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l291_c11_0a6c]
signal BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l291_c7_c678]
signal n8_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l291_c7_c678]
signal t8_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l291_c7_c678]
signal result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l291_c7_c678]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l291_c7_c678]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l291_c7_c678]
signal result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l291_c7_c678]
signal result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l291_c7_c678]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l294_c11_f14a]
signal BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l294_c7_7ea5]
signal n8_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l294_c7_7ea5]
signal t8_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l294_c7_7ea5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l294_c7_7ea5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l294_c7_7ea5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l294_c7_7ea5]
signal result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l294_c7_7ea5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l294_c7_7ea5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l297_c30_4ec1]
signal sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l302_c11_4c90]
signal BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l302_c7_69b8]
signal n8_MUX_uxn_opcodes_h_l302_c7_69b8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l302_c7_69b8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l302_c7_69b8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l302_c7_69b8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l302_c7_69b8]
signal result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l302_c7_69b8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l302_c7_69b8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l308_c11_5332]
signal BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l308_c7_846f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l308_c7_846f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l308_c7_846f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l308_c7_846f]
signal result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l312_c11_5064]
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l312_c7_3b23]
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l312_c7_3b23]
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c551( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf
BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_left,
BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_right,
BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_return_output);

-- n8_MUX_uxn_opcodes_h_l286_c2_7f12
n8_MUX_uxn_opcodes_h_l286_c2_7f12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l286_c2_7f12_cond,
n8_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue,
n8_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse,
n8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output);

-- t8_MUX_uxn_opcodes_h_l286_c2_7f12
t8_MUX_uxn_opcodes_h_l286_c2_7f12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l286_c2_7f12_cond,
t8_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue,
t8_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse,
t8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12
result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12
result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12
result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_cond,
result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12
result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12
result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output);

-- printf_uxn_opcodes_h_l287_c3_ed90_uxn_opcodes_h_l287_c3_ed90
printf_uxn_opcodes_h_l287_c3_ed90_uxn_opcodes_h_l287_c3_ed90 : entity work.printf_uxn_opcodes_h_l287_c3_ed90_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l287_c3_ed90_uxn_opcodes_h_l287_c3_ed90_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c
BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_left,
BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_right,
BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output);

-- n8_MUX_uxn_opcodes_h_l291_c7_c678
n8_MUX_uxn_opcodes_h_l291_c7_c678 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l291_c7_c678_cond,
n8_MUX_uxn_opcodes_h_l291_c7_c678_iftrue,
n8_MUX_uxn_opcodes_h_l291_c7_c678_iffalse,
n8_MUX_uxn_opcodes_h_l291_c7_c678_return_output);

-- t8_MUX_uxn_opcodes_h_l291_c7_c678
t8_MUX_uxn_opcodes_h_l291_c7_c678 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l291_c7_c678_cond,
t8_MUX_uxn_opcodes_h_l291_c7_c678_iftrue,
t8_MUX_uxn_opcodes_h_l291_c7_c678_iffalse,
t8_MUX_uxn_opcodes_h_l291_c7_c678_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678
result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678
result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678
result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_cond,
result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678
result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678
result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a
BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_left,
BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_right,
BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output);

-- n8_MUX_uxn_opcodes_h_l294_c7_7ea5
n8_MUX_uxn_opcodes_h_l294_c7_7ea5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l294_c7_7ea5_cond,
n8_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue,
n8_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse,
n8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output);

-- t8_MUX_uxn_opcodes_h_l294_c7_7ea5
t8_MUX_uxn_opcodes_h_l294_c7_7ea5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l294_c7_7ea5_cond,
t8_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue,
t8_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse,
t8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5
result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5
result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5
result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_cond,
result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5
result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5
result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output);

-- sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1
sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_ins,
sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_x,
sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_y,
sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90
BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_left,
BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_right,
BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_return_output);

-- n8_MUX_uxn_opcodes_h_l302_c7_69b8
n8_MUX_uxn_opcodes_h_l302_c7_69b8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l302_c7_69b8_cond,
n8_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue,
n8_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse,
n8_MUX_uxn_opcodes_h_l302_c7_69b8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8
result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8
result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_cond,
result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8
result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8
result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332
BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_left,
BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_right,
BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f
result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f
result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f
result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_cond,
result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064
BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_left,
BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_right,
BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_return_output,
 n8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output,
 t8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output,
 n8_MUX_uxn_opcodes_h_l291_c7_c678_return_output,
 t8_MUX_uxn_opcodes_h_l291_c7_c678_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output,
 n8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output,
 t8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output,
 sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_return_output,
 n8_MUX_uxn_opcodes_h_l302_c7_69b8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l288_c3_936e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l287_c3_ed90_uxn_opcodes_h_l287_c3_ed90_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l292_c3_f861 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l302_c7_69b8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l299_c3_76b0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l302_c7_69b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l305_c3_b27f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_d54f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l308_c7_846f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l312_l308_l302_l291_l286_DUPLICATE_365f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l291_l294_l286_DUPLICATE_0b0d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l291_l308_l286_DUPLICATE_6c39_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l302_l291_l286_DUPLICATE_7483_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l312_l308_l302_l294_l291_DUPLICATE_8d76_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l317_l282_DUPLICATE_febb_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l288_c3_936e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l288_c3_936e;
     VAR_sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l292_c3_f861 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l292_c3_f861;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l305_c3_b27f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l305_c3_b27f;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l299_c3_76b0 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l299_c3_76b0;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_d54f := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_d54f;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l291_c7_c678_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse := n8;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l291_c7_c678_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l297_c30_4ec1] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_ins;
     sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_x <= VAR_sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_x;
     sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_y <= VAR_sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_return_output := sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l308_c7_846f] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l308_c7_846f_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l302_c11_4c90] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_left;
     BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_return_output := BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l312_c11_5064] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_left;
     BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_return_output := BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l312_l308_l302_l291_l286_DUPLICATE_365f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l312_l308_l302_l291_l286_DUPLICATE_365f_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l302_l291_l286_DUPLICATE_7483 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l302_l291_l286_DUPLICATE_7483_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l286_c6_85cf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_left;
     BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output := BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l291_l308_l286_DUPLICATE_6c39 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l291_l308_l286_DUPLICATE_6c39_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l291_c11_0a6c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_left;
     BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output := BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l312_l308_l302_l294_l291_DUPLICATE_8d76 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l312_l308_l302_l294_l291_DUPLICATE_8d76_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l291_l294_l286_DUPLICATE_0b0d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l291_l294_l286_DUPLICATE_0b0d_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l294_c11_f14a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_left;
     BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output := BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l308_c11_5332] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_left;
     BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_return_output := BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l286_c2_7f12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l286_c2_7f12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l286_c6_85cf_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l291_c7_c678_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l291_c7_c678_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l291_c11_0a6c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l294_c7_7ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l294_c7_7ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l294_c11_f14a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l302_c7_69b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c11_4c90_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l308_c11_5332_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_5064_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l291_l294_l286_DUPLICATE_0b0d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l291_l294_l286_DUPLICATE_0b0d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l291_l294_l286_DUPLICATE_0b0d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l312_l308_l302_l294_l291_DUPLICATE_8d76_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l312_l308_l302_l294_l291_DUPLICATE_8d76_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l312_l308_l302_l294_l291_DUPLICATE_8d76_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l312_l308_l302_l294_l291_DUPLICATE_8d76_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l312_l308_l302_l294_l291_DUPLICATE_8d76_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l302_l291_l286_DUPLICATE_7483_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l302_l291_l286_DUPLICATE_7483_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l302_l291_l286_DUPLICATE_7483_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l312_l308_l302_l291_l286_DUPLICATE_365f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l312_l308_l302_l291_l286_DUPLICATE_365f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l312_l308_l302_l291_l286_DUPLICATE_365f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l312_l308_l302_l291_l286_DUPLICATE_365f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l312_l308_l302_l291_l286_DUPLICATE_365f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l291_l308_l286_DUPLICATE_6c39_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l291_l308_l286_DUPLICATE_6c39_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l291_l308_l286_DUPLICATE_6c39_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l308_c7_846f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l297_c30_4ec1_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l312_c7_3b23] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_return_output;

     -- n8_MUX[uxn_opcodes_h_l302_c7_69b8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l302_c7_69b8_cond <= VAR_n8_MUX_uxn_opcodes_h_l302_c7_69b8_cond;
     n8_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue;
     n8_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l302_c7_69b8_return_output := n8_MUX_uxn_opcodes_h_l302_c7_69b8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l308_c7_846f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_return_output := result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l302_c7_69b8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l308_c7_846f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_return_output;

     -- t8_MUX[uxn_opcodes_h_l294_c7_7ea5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l294_c7_7ea5_cond <= VAR_t8_MUX_uxn_opcodes_h_l294_c7_7ea5_cond;
     t8_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue;
     t8_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output := t8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l286_c1_1890] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l294_c7_7ea5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l312_c7_3b23] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l287_c3_ed90_uxn_opcodes_h_l287_c3_ed90_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l286_c1_1890_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l302_c7_69b8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_3b23_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l302_c7_69b8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_3b23_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l308_c7_846f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l308_c7_846f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l291_c7_c678_iffalse := VAR_t8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;
     -- printf_uxn_opcodes_h_l287_c3_ed90[uxn_opcodes_h_l287_c3_ed90] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l287_c3_ed90_uxn_opcodes_h_l287_c3_ed90_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l287_c3_ed90_uxn_opcodes_h_l287_c3_ed90_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- t8_MUX[uxn_opcodes_h_l291_c7_c678] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l291_c7_c678_cond <= VAR_t8_MUX_uxn_opcodes_h_l291_c7_c678_cond;
     t8_MUX_uxn_opcodes_h_l291_c7_c678_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l291_c7_c678_iftrue;
     t8_MUX_uxn_opcodes_h_l291_c7_c678_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l291_c7_c678_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l291_c7_c678_return_output := t8_MUX_uxn_opcodes_h_l291_c7_c678_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l291_c7_c678] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output;

     -- n8_MUX[uxn_opcodes_h_l294_c7_7ea5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l294_c7_7ea5_cond <= VAR_n8_MUX_uxn_opcodes_h_l294_c7_7ea5_cond;
     n8_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue;
     n8_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output := n8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l294_c7_7ea5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l302_c7_69b8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_return_output := result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l308_c7_846f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l308_c7_846f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l302_c7_69b8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l291_c7_c678_iffalse := VAR_n8_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l308_c7_846f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l308_c7_846f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c7_69b8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c7_69b8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse := VAR_t8_MUX_uxn_opcodes_h_l291_c7_c678_return_output;
     -- t8_MUX[uxn_opcodes_h_l286_c2_7f12] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l286_c2_7f12_cond <= VAR_t8_MUX_uxn_opcodes_h_l286_c2_7f12_cond;
     t8_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue;
     t8_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output := t8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l294_c7_7ea5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;

     -- n8_MUX[uxn_opcodes_h_l291_c7_c678] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l291_c7_c678_cond <= VAR_n8_MUX_uxn_opcodes_h_l291_c7_c678_cond;
     n8_MUX_uxn_opcodes_h_l291_c7_c678_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l291_c7_c678_iftrue;
     n8_MUX_uxn_opcodes_h_l291_c7_c678_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l291_c7_c678_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l291_c7_c678_return_output := n8_MUX_uxn_opcodes_h_l291_c7_c678_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l302_c7_69b8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l302_c7_69b8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l294_c7_7ea5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output := result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l291_c7_c678] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l286_c2_7f12] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse := VAR_n8_MUX_uxn_opcodes_h_l291_c7_c678_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c7_69b8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l291_c7_c678_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c7_69b8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output;
     -- n8_MUX[uxn_opcodes_h_l286_c2_7f12] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l286_c2_7f12_cond <= VAR_n8_MUX_uxn_opcodes_h_l286_c2_7f12_cond;
     n8_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue;
     n8_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output := n8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l291_c7_c678] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_cond;
     result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_return_output := result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l286_c2_7f12] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l294_c7_7ea5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l291_c7_c678] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l294_c7_7ea5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l286_c2_7f12_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l294_c7_7ea5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l291_c7_c678_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l291_c7_c678_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l291_c7_c678] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l291_c7_c678] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l286_c2_7f12] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_cond;
     result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_return_output := result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l286_c2_7f12] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l291_c7_c678_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l291_c7_c678_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l286_c2_7f12] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l286_c2_7f12] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l317_l282_DUPLICATE_febb LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l317_l282_DUPLICATE_febb_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c551(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l286_c2_7f12_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l286_c2_7f12_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l286_c2_7f12_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l286_c2_7f12_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l286_c2_7f12_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l317_l282_DUPLICATE_febb_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l317_l282_DUPLICATE_febb_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
