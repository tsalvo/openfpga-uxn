-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 79
entity eor2_0CLK_f74041be is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor2_0CLK_f74041be;
architecture arch of eor2_0CLK_f74041be is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1067_c6_3694]
signal BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1067_c1_3ac8]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1067_c2_408b]
signal tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1067_c2_408b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1067_c2_408b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1067_c2_408b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1067_c2_408b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1067_c2_408b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1067_c2_408b]
signal result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l1067_c2_408b]
signal t16_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(15 downto 0);

-- n16_MUX[uxn_opcodes_h_l1067_c2_408b]
signal n16_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l1068_c3_7fb3[uxn_opcodes_h_l1068_c3_7fb3]
signal printf_uxn_opcodes_h_l1068_c3_7fb3_uxn_opcodes_h_l1068_c3_7fb3_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1072_c11_2889]
signal BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1072_c7_f1e3]
signal tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1072_c7_f1e3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1072_c7_f1e3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1072_c7_f1e3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1072_c7_f1e3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1072_c7_f1e3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1072_c7_f1e3]
signal result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l1072_c7_f1e3]
signal t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(15 downto 0);

-- n16_MUX[uxn_opcodes_h_l1072_c7_f1e3]
signal n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1075_c11_1b58]
signal BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1075_c7_98e3]
signal tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1075_c7_98e3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1075_c7_98e3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1075_c7_98e3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1075_c7_98e3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1075_c7_98e3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1075_c7_98e3]
signal result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l1075_c7_98e3]
signal t16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(15 downto 0);

-- n16_MUX[uxn_opcodes_h_l1075_c7_98e3]
signal n16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1080_c11_d07f]
signal BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1080_c7_dfd4]
signal tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1080_c7_dfd4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1080_c7_dfd4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1080_c7_dfd4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1080_c7_dfd4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1080_c7_dfd4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1080_c7_dfd4]
signal result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l1080_c7_dfd4]
signal t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(15 downto 0);

-- n16_MUX[uxn_opcodes_h_l1080_c7_dfd4]
signal n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l1081_c3_f1ca]
signal BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1084_c11_23e7]
signal BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1084_c7_84e2]
signal tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1084_c7_84e2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1084_c7_84e2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1084_c7_84e2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1084_c7_84e2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1084_c7_84e2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1084_c7_84e2]
signal result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(7 downto 0);

-- n16_MUX[uxn_opcodes_h_l1084_c7_84e2]
signal n16_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1088_c11_8d66]
signal BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1088_c7_9cdc]
signal tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1088_c7_9cdc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1088_c7_9cdc]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1088_c7_9cdc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1088_c7_9cdc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1088_c7_9cdc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1088_c7_9cdc]
signal result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(7 downto 0);

-- n16_MUX[uxn_opcodes_h_l1088_c7_9cdc]
signal n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l1089_c3_24a3]
signal BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_return_output : unsigned(15 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1090_c11_55e3]
signal BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_left : unsigned(15 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_right : unsigned(15 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1092_c30_6faf]
signal sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1097_c11_3d37]
signal BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1097_c7_6983]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1097_c7_6983]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1097_c7_6983]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1097_c7_6983]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1097_c7_6983]
signal result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_return_output : unsigned(7 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l1100_c31_ff18]
signal CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1102_c11_0425]
signal BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1102_c7_babc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1102_c7_babc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_return_output : unsigned(0 downto 0);

-- CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2
signal CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_x : unsigned(15 downto 0);
signal CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_return_output : unsigned(15 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_8c29( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694
BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_left,
BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_right,
BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1067_c2_408b
tmp16_MUX_uxn_opcodes_h_l1067_c2_408b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_cond,
tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue,
tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse,
tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b
result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b
result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_return_output);

-- t16_MUX_uxn_opcodes_h_l1067_c2_408b
t16_MUX_uxn_opcodes_h_l1067_c2_408b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1067_c2_408b_cond,
t16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue,
t16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse,
t16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output);

-- n16_MUX_uxn_opcodes_h_l1067_c2_408b
n16_MUX_uxn_opcodes_h_l1067_c2_408b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1067_c2_408b_cond,
n16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue,
n16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse,
n16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output);

-- printf_uxn_opcodes_h_l1068_c3_7fb3_uxn_opcodes_h_l1068_c3_7fb3
printf_uxn_opcodes_h_l1068_c3_7fb3_uxn_opcodes_h_l1068_c3_7fb3 : entity work.printf_uxn_opcodes_h_l1068_c3_7fb3_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1068_c3_7fb3_uxn_opcodes_h_l1068_c3_7fb3_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889
BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_left,
BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_right,
BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3
tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond,
tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue,
tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse,
tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3
result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3
result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3
result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3
result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3
result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond,
result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output);

-- t16_MUX_uxn_opcodes_h_l1072_c7_f1e3
t16_MUX_uxn_opcodes_h_l1072_c7_f1e3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond,
t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue,
t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse,
t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output);

-- n16_MUX_uxn_opcodes_h_l1072_c7_f1e3
n16_MUX_uxn_opcodes_h_l1072_c7_f1e3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond,
n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue,
n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse,
n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58
BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_left,
BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_right,
BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3
tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond,
tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue,
tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse,
tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3
result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3
result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3
result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3
result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3
result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_cond,
result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output);

-- t16_MUX_uxn_opcodes_h_l1075_c7_98e3
t16_MUX_uxn_opcodes_h_l1075_c7_98e3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond,
t16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue,
t16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse,
t16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output);

-- n16_MUX_uxn_opcodes_h_l1075_c7_98e3
n16_MUX_uxn_opcodes_h_l1075_c7_98e3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond,
n16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue,
n16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse,
n16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f
BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_left,
BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_right,
BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4
tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond,
tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue,
tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse,
tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4
result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4
result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4
result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4
result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output);

-- t16_MUX_uxn_opcodes_h_l1080_c7_dfd4
t16_MUX_uxn_opcodes_h_l1080_c7_dfd4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond,
t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue,
t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse,
t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output);

-- n16_MUX_uxn_opcodes_h_l1080_c7_dfd4
n16_MUX_uxn_opcodes_h_l1080_c7_dfd4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond,
n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue,
n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse,
n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca
BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_left,
BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_right,
BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7
BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_left,
BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_right,
BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2
tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_cond,
tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue,
tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse,
tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2
result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2
result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2
result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2
result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output);

-- n16_MUX_uxn_opcodes_h_l1084_c7_84e2
n16_MUX_uxn_opcodes_h_l1084_c7_84e2 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1084_c7_84e2_cond,
n16_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue,
n16_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse,
n16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66
BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_left,
BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_right,
BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc
tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond,
tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue,
tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse,
tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc
result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc
result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc
result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc
result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc
result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond,
result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output);

-- n16_MUX_uxn_opcodes_h_l1088_c7_9cdc
n16_MUX_uxn_opcodes_h_l1088_c7_9cdc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond,
n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue,
n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse,
n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3
BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_left,
BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_right,
BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3
BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3 : entity work.BIN_OP_XOR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_left,
BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_right,
BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf
sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_ins,
sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_x,
sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_y,
sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37
BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_left,
BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_right,
BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983
result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983
result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983
result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983
result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_cond,
result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_return_output);

-- CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18
CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18_x,
CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425
BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_left,
BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_right,
BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc
result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc
result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_return_output);

-- CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2
CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_x,
CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_return_output,
 tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
 t16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
 n16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output,
 tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output,
 t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output,
 n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output,
 tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output,
 t16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output,
 n16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output,
 tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output,
 t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output,
 n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output,
 BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output,
 tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output,
 n16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output,
 tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output,
 n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output,
 BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_return_output,
 sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_return_output,
 CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_return_output,
 CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_iffalse : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1069_c3_6616 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1067_c2_408b_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1068_c3_7fb3_uxn_opcodes_h_l1068_c3_7fb3_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1073_c3_3c25 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1078_c3_13ba : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1082_c3_0c9c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1084_c7_84e2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1094_c3_67da : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_return_output : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1095_c21_7f0a_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1099_c3_a6b5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1100_c21_a1c2_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_a228_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1072_l1102_l1067_l1097_l1084_l1080_l1075_DUPLICATE_4f2d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1072_l1067_l1088_l1084_l1080_l1075_DUPLICATE_e865_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_190f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1072_l1102_l1097_l1088_l1084_l1080_l1075_DUPLICATE_b404_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1081_l1089_l1076_l1085_DUPLICATE_f14d_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_x : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1097_l1084_DUPLICATE_4682_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1107_l1063_DUPLICATE_c2ca_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1073_c3_3c25 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1073_c3_3c25;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1082_c3_0c9c := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1082_c3_0c9c;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1094_c3_67da := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1094_c3_67da;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1078_c3_13ba := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1078_c3_13ba;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1099_c3_a6b5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1099_c3_a6b5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_right := to_unsigned(6, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1069_c3_6616 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1069_c3_6616;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_right := to_unsigned(7, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_ins := VAR_ins;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_left := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_left := t16;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_right := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse := t16;
     VAR_CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18_x := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse := tmp16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_a228 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_a228_return_output := result.is_sp_shift;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1081_l1089_l1076_l1085_DUPLICATE_f14d LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1081_l1089_l1076_l1085_DUPLICATE_f14d_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1075_c11_1b58] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_left;
     BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output := BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1072_l1102_l1067_l1097_l1084_l1080_l1075_DUPLICATE_4f2d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1072_l1102_l1067_l1097_l1084_l1080_l1075_DUPLICATE_4f2d_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1097_c11_3d37] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_left;
     BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_return_output := BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1097_l1084_DUPLICATE_4682 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1097_l1084_DUPLICATE_4682_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1072_l1067_l1088_l1084_l1080_l1075_DUPLICATE_e865 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1072_l1067_l1088_l1084_l1080_l1075_DUPLICATE_e865_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l1092_c30_6faf] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_ins;
     sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_x;
     sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_return_output := sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1080_c11_d07f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output;

     -- CONST_SR_8[uxn_opcodes_h_l1100_c31_ff18] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18_x <= VAR_CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18_return_output := CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1084_c11_23e7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_left;
     BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output := BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1102_c11_0425] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_left;
     BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_return_output := BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1088_c11_8d66] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_left;
     BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output := BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1067_c6_3694] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_left;
     BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output := BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1072_c11_2889] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_left;
     BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output := BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_190f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_190f_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1072_l1102_l1097_l1088_l1084_l1080_l1075_DUPLICATE_b404 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1072_l1102_l1097_l1088_l1084_l1080_l1075_DUPLICATE_b404_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1067_c2_408b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1067_c2_408b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c6_3694_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1072_c11_2889_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1075_c11_1b58_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1080_c11_d07f_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1084_c7_84e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1084_c11_23e7_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1088_c11_8d66_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1097_c11_3d37_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1102_c11_0425_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1081_l1089_l1076_l1085_DUPLICATE_f14d_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1081_l1089_l1076_l1085_DUPLICATE_f14d_return_output;
     VAR_CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1081_l1089_l1076_l1085_DUPLICATE_f14d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1072_l1067_l1088_l1084_l1080_l1075_DUPLICATE_e865_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1072_l1067_l1088_l1084_l1080_l1075_DUPLICATE_e865_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1072_l1067_l1088_l1084_l1080_l1075_DUPLICATE_e865_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1072_l1067_l1088_l1084_l1080_l1075_DUPLICATE_e865_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1072_l1067_l1088_l1084_l1080_l1075_DUPLICATE_e865_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1072_l1067_l1088_l1084_l1080_l1075_DUPLICATE_e865_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1072_l1102_l1097_l1088_l1084_l1080_l1075_DUPLICATE_b404_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1072_l1102_l1097_l1088_l1084_l1080_l1075_DUPLICATE_b404_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1072_l1102_l1097_l1088_l1084_l1080_l1075_DUPLICATE_b404_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1072_l1102_l1097_l1088_l1084_l1080_l1075_DUPLICATE_b404_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1072_l1102_l1097_l1088_l1084_l1080_l1075_DUPLICATE_b404_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1072_l1102_l1097_l1088_l1084_l1080_l1075_DUPLICATE_b404_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1072_l1102_l1097_l1088_l1084_l1080_l1075_DUPLICATE_b404_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_a228_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_a228_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_a228_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_a228_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_a228_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_a228_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1072_l1102_l1067_l1097_l1084_l1080_l1075_DUPLICATE_4f2d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1072_l1102_l1067_l1097_l1084_l1080_l1075_DUPLICATE_4f2d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1072_l1102_l1067_l1097_l1084_l1080_l1075_DUPLICATE_4f2d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1072_l1102_l1067_l1097_l1084_l1080_l1075_DUPLICATE_4f2d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1072_l1102_l1067_l1097_l1084_l1080_l1075_DUPLICATE_4f2d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1072_l1102_l1067_l1097_l1084_l1080_l1075_DUPLICATE_4f2d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1072_l1102_l1067_l1097_l1084_l1080_l1075_DUPLICATE_4f2d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1097_l1084_DUPLICATE_4682_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1097_l1084_DUPLICATE_4682_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_190f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_190f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_190f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_190f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_190f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1072_l1067_l1097_l1084_l1080_l1075_DUPLICATE_190f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1092_c30_6faf_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1097_c7_6983] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1088_c7_9cdc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1067_c1_3ac8] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1102_c7_babc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_return_output;

     -- CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2 LATENCY=0
     -- Inputs
     CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_x <= VAR_CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_x;
     -- Outputs
     VAR_CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_return_output := CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l1100_c21_a1c2] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1100_c21_a1c2_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l1100_c31_ff18_return_output);

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1102_c7_babc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1097_c7_6983] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l1089_c3_24a3] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_left;
     BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_return_output := BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l1081_c3_f1ca] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_left;
     BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_return_output := BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l1081_c3_f1ca_return_output;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_left := VAR_BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l1089_c3_24a3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1100_c21_a1c2_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue := VAR_CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue := VAR_CONST_SL_8_uint16_t_uxn_opcodes_h_l1077_l1086_DUPLICATE_0ea2_return_output;
     VAR_printf_uxn_opcodes_h_l1068_c3_7fb3_uxn_opcodes_h_l1068_c3_7fb3_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1067_c1_3ac8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1102_c7_babc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1097_c7_6983_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1102_c7_babc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1097_c7_6983_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1088_c7_9cdc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1097_c7_6983] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_return_output;

     -- t16_MUX[uxn_opcodes_h_l1080_c7_dfd4] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond <= VAR_t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond;
     t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue;
     t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output := t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1088_c7_9cdc] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;

     -- BIN_OP_XOR[uxn_opcodes_h_l1090_c11_55e3] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_left;
     BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_return_output := BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1097_c7_6983] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_return_output := result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1084_c7_84e2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;

     -- printf_uxn_opcodes_h_l1068_c3_7fb3[uxn_opcodes_h_l1068_c3_7fb3] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1068_c3_7fb3_uxn_opcodes_h_l1068_c3_7fb3_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1068_c3_7fb3_uxn_opcodes_h_l1068_c3_7fb3_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- n16_MUX[uxn_opcodes_h_l1088_c7_9cdc] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond <= VAR_n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond;
     n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue;
     n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output := n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1097_c7_6983] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_return_output;

     -- Submodule level 3
     VAR_tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1097_c7_6983_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1097_c7_6983_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1097_c7_6983_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;
     -- n16_MUX[uxn_opcodes_h_l1084_c7_84e2] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1084_c7_84e2_cond <= VAR_n16_MUX_uxn_opcodes_h_l1084_c7_84e2_cond;
     n16_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue;
     n16_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output := n16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1088_c7_9cdc] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond;
     tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output := tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;

     -- t16_MUX[uxn_opcodes_h_l1075_c7_98e3] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond <= VAR_t16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond;
     t16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue;
     t16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output := t16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1084_c7_84e2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1088_c7_9cdc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1084_c7_84e2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l1095_c21_7f0a] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1095_c21_7f0a_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1090_c11_55e3_return_output);

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1088_c7_9cdc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1080_c7_dfd4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;

     -- Submodule level 4
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1095_c21_7f0a_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1088_c7_9cdc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output := result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;

     -- n16_MUX[uxn_opcodes_h_l1080_c7_dfd4] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond <= VAR_n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond;
     n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue;
     n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output := n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1084_c7_84e2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1075_c7_98e3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1080_c7_dfd4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;

     -- t16_MUX[uxn_opcodes_h_l1072_c7_f1e3] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond <= VAR_t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond;
     t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue;
     t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output := t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1080_c7_dfd4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1084_c7_84e2] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_cond;
     tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output := tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1084_c7_84e2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;

     -- Submodule level 5
     VAR_n16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1088_c7_9cdc_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1072_c7_f1e3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;

     -- n16_MUX[uxn_opcodes_h_l1075_c7_98e3] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond <= VAR_n16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond;
     n16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue;
     n16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output := n16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1080_c7_dfd4] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond;
     tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output := tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;

     -- t16_MUX[uxn_opcodes_h_l1067_c2_408b] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1067_c2_408b_cond <= VAR_t16_MUX_uxn_opcodes_h_l1067_c2_408b_cond;
     t16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue;
     t16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output := t16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1075_c7_98e3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1075_c7_98e3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1084_c7_84e2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1080_c7_dfd4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1080_c7_dfd4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;

     -- Submodule level 6
     VAR_n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1084_c7_84e2_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1067_c2_408b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1080_c7_dfd4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1072_c7_f1e3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1075_c7_98e3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;

     -- n16_MUX[uxn_opcodes_h_l1072_c7_f1e3] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond <= VAR_n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond;
     n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue;
     n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output := n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1075_c7_98e3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1075_c7_98e3] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_cond;
     tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output := tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1072_c7_f1e3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;

     -- Submodule level 7
     VAR_n16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1080_c7_dfd4_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l1072_c7_f1e3] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond;
     tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output := tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1075_c7_98e3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output := result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1067_c2_408b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_return_output;

     -- n16_MUX[uxn_opcodes_h_l1067_c2_408b] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1067_c2_408b_cond <= VAR_n16_MUX_uxn_opcodes_h_l1067_c2_408b_cond;
     n16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue;
     n16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output := n16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1072_c7_f1e3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1072_c7_f1e3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1067_c2_408b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output;

     -- Submodule level 8
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1075_c7_98e3_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l1067_c2_408b] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_cond;
     tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output := tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1067_c2_408b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1067_c2_408b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1072_c7_f1e3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output := result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;

     -- Submodule level 9
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1072_c7_f1e3_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l1067_c2_408b_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1067_c2_408b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_return_output;

     -- Submodule level 10
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1107_l1063_DUPLICATE_c2ca LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1107_l1063_DUPLICATE_c2ca_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8c29(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c2_408b_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1067_c2_408b_return_output);

     -- Submodule level 11
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1107_l1063_DUPLICATE_c2ca_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1107_l1063_DUPLICATE_c2ca_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
