-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 55
entity sth_0CLK_edc09f97 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth_0CLK_edc09f97;
architecture arch of sth_0CLK_edc09f97 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2729_c6_b199]
signal BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2729_c1_cf07]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2729_c2_ea1b]
signal t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2729_c2_ea1b]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2729_c2_ea1b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2729_c2_ea1b]
signal result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2729_c2_ea1b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2729_c2_ea1b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2729_c2_ea1b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2729_c2_ea1b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2729_c2_ea1b]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l2730_c3_5f91[uxn_opcodes_h_l2730_c3_5f91]
signal printf_uxn_opcodes_h_l2730_c3_5f91_uxn_opcodes_h_l2730_c3_5f91_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2735_c11_5590]
signal BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2735_c7_652c]
signal t8_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2735_c7_652c]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2735_c7_652c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2735_c7_652c]
signal result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2735_c7_652c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2735_c7_652c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2735_c7_652c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2735_c7_652c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2735_c7_652c]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2738_c11_e9b0]
signal BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2738_c7_1f6e]
signal t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2738_c7_1f6e]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2738_c7_1f6e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2738_c7_1f6e]
signal result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2738_c7_1f6e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2738_c7_1f6e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2738_c7_1f6e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2738_c7_1f6e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2738_c7_1f6e]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2742_c32_86c6]
signal BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l2742_c32_e20d]
signal BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l2742_c32_63d3]
signal MUX_uxn_opcodes_h_l2742_c32_63d3_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2742_c32_63d3_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2742_c32_63d3_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2742_c32_63d3_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2744_c11_2a7f]
signal BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2744_c7_3775]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : signed(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2744_c7_3775]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2744_c7_3775]
signal result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2744_c7_3775]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2744_c7_3775]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2744_c7_3775]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2744_c7_3775]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2748_c11_c0de]
signal BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2748_c7_e6b6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2748_c7_e6b6]
signal result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2748_c7_e6b6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2748_c7_e6b6]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2748_c7_e6b6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2748_c7_e6b6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2754_c11_7d63]
signal BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2754_c7_0dfe]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2754_c7_0dfe]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2754_c7_0dfe]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_f6cd( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : signed;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_read := ref_toks_1;
      base.sp_relative_shift := ref_toks_2;
      base.stack_value := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_stack_write := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199
BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_left,
BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_right,
BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_return_output);

-- t8_MUX_uxn_opcodes_h_l2729_c2_ea1b
t8_MUX_uxn_opcodes_h_l2729_c2_ea1b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond,
t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue,
t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse,
t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b
result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b
result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond,
result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b
result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b
result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b
result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output);

-- printf_uxn_opcodes_h_l2730_c3_5f91_uxn_opcodes_h_l2730_c3_5f91
printf_uxn_opcodes_h_l2730_c3_5f91_uxn_opcodes_h_l2730_c3_5f91 : entity work.printf_uxn_opcodes_h_l2730_c3_5f91_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2730_c3_5f91_uxn_opcodes_h_l2730_c3_5f91_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590
BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_left,
BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_right,
BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output);

-- t8_MUX_uxn_opcodes_h_l2735_c7_652c
t8_MUX_uxn_opcodes_h_l2735_c7_652c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2735_c7_652c_cond,
t8_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue,
t8_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse,
t8_MUX_uxn_opcodes_h_l2735_c7_652c_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c
result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c
result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_cond,
result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c
result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c
result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c
result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_left,
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_right,
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output);

-- t8_MUX_uxn_opcodes_h_l2738_c7_1f6e
t8_MUX_uxn_opcodes_h_l2738_c7_1f6e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond,
t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue,
t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse,
t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e
result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e
result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond,
result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e
result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6
BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_left,
BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_right,
BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d
BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_left,
BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_right,
BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_return_output);

-- MUX_uxn_opcodes_h_l2742_c32_63d3
MUX_uxn_opcodes_h_l2742_c32_63d3 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2742_c32_63d3_cond,
MUX_uxn_opcodes_h_l2742_c32_63d3_iftrue,
MUX_uxn_opcodes_h_l2742_c32_63d3_iffalse,
MUX_uxn_opcodes_h_l2742_c32_63d3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f
BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_left,
BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_right,
BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775
result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775
result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775
result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_cond,
result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775
result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775
result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de
BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_left,
BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_right,
BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6
result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6
result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond,
result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6
result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6
result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63
BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_left,
BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_right,
BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe
result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe
result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_return_output,
 t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output,
 t8_MUX_uxn_opcodes_h_l2735_c7_652c_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output,
 t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_return_output,
 BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_return_output,
 MUX_uxn_opcodes_h_l2742_c32_63d3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2732_c3_c011 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2730_c3_5f91_uxn_opcodes_h_l2730_c3_5f91_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2736_c3_e91a : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2742_c32_63d3_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2742_c32_63d3_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2742_c32_63d3_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2742_c32_63d3_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2746_c3_6b32 : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2751_c3_7eb3 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2735_l2729_l2744_DUPLICATE_7150_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2729_DUPLICATE_de0f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2735_l2748_l2729_l2744_DUPLICATE_e103_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2744_l2738_l2735_l2729_l2754_DUPLICATE_8386_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2748_l2738_l2735_l2729_l2754_DUPLICATE_5228_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2735_l2738_DUPLICATE_5b3e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2754_DUPLICATE_cdc6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2748_l2738_l2744_DUPLICATE_3bac_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f6cd_uxn_opcodes_h_l2760_l2725_DUPLICATE_924a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l2742_c32_63d3_iffalse := resize(to_signed(-1, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2751_c3_7eb3 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2751_c3_7eb3;
     VAR_BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_right := to_unsigned(5, 3);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2746_c3_6b32 := signed(std_logic_vector(resize(to_unsigned(2, 2), 8)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2746_c3_6b32;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2736_c3_e91a := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2736_c3_e91a;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2732_c3_c011 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2732_c3_c011;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_right := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l2742_c32_63d3_iftrue := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_right := to_unsigned(1, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_right := to_unsigned(128, 8);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2754_DUPLICATE_cdc6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2754_DUPLICATE_cdc6_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2748_l2738_l2735_l2729_l2754_DUPLICATE_5228 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2748_l2738_l2735_l2729_l2754_DUPLICATE_5228_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2735_l2748_l2729_l2744_DUPLICATE_e103 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2735_l2748_l2729_l2744_DUPLICATE_e103_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2735_c11_5590] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_left;
     BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output := BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2744_c11_2a7f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2738_c11_e9b0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2748_c11_c0de] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_left;
     BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_return_output := BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2748_l2738_l2744_DUPLICATE_3bac LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2748_l2738_l2744_DUPLICATE_3bac_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2729_c6_b199] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_left;
     BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output := BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2729_DUPLICATE_de0f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2729_DUPLICATE_de0f_return_output := result.stack_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2735_l2738_DUPLICATE_5b3e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2735_l2738_DUPLICATE_5b3e_return_output := result.is_stack_read;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2744_l2738_l2735_l2729_l2754_DUPLICATE_8386 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2744_l2738_l2735_l2729_l2754_DUPLICATE_8386_return_output := result.is_stack_write;

     -- BIN_OP_AND[uxn_opcodes_h_l2742_c32_86c6] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_left;
     BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_return_output := BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2754_c11_7d63] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_left;
     BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_return_output := BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2735_l2729_l2744_DUPLICATE_7150 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2735_l2729_l2744_DUPLICATE_7150_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_left := VAR_BIN_OP_AND_uxn_opcodes_h_l2742_c32_86c6_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2729_c6_b199_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2735_c7_652c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2735_c11_5590_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_e9b0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2744_c11_2a7f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2748_c11_c0de_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2754_c11_7d63_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2735_l2729_l2744_DUPLICATE_7150_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2735_l2729_l2744_DUPLICATE_7150_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2735_l2729_l2744_DUPLICATE_7150_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2754_DUPLICATE_cdc6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2754_DUPLICATE_cdc6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2754_DUPLICATE_cdc6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2754_DUPLICATE_cdc6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2754_DUPLICATE_cdc6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2735_l2748_l2729_l2744_DUPLICATE_e103_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2735_l2748_l2729_l2744_DUPLICATE_e103_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2735_l2748_l2729_l2744_DUPLICATE_e103_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2735_l2748_l2729_l2744_DUPLICATE_e103_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2748_l2738_l2735_l2729_l2754_DUPLICATE_5228_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2748_l2738_l2735_l2729_l2754_DUPLICATE_5228_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2748_l2738_l2735_l2729_l2754_DUPLICATE_5228_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2748_l2738_l2735_l2729_l2754_DUPLICATE_5228_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2748_l2738_l2735_l2729_l2754_DUPLICATE_5228_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2735_l2738_DUPLICATE_5b3e_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2735_l2738_DUPLICATE_5b3e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2744_l2738_l2735_l2729_l2754_DUPLICATE_8386_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2744_l2738_l2735_l2729_l2754_DUPLICATE_8386_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2744_l2738_l2735_l2729_l2754_DUPLICATE_8386_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2744_l2738_l2735_l2729_l2754_DUPLICATE_8386_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2744_l2738_l2735_l2729_l2754_DUPLICATE_8386_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2748_l2738_l2744_DUPLICATE_3bac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2748_l2738_l2744_DUPLICATE_3bac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2748_l2738_l2744_DUPLICATE_3bac_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2729_DUPLICATE_de0f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2729_DUPLICATE_de0f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2729_DUPLICATE_de0f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2729_DUPLICATE_de0f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2748_l2744_l2738_l2735_l2729_DUPLICATE_de0f_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2754_c7_0dfe] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2754_c7_0dfe] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output;

     -- t8_MUX[uxn_opcodes_h_l2738_c7_1f6e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond <= VAR_t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond;
     t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue;
     t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output := t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2729_c1_cf07] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2748_c7_e6b6] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output := result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l2742_c32_e20d] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_left;
     BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_return_output := BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2744_c7_3775] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2748_c7_e6b6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2738_c7_1f6e] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2748_c7_e6b6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2754_c7_0dfe] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l2742_c32_63d3_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l2742_c32_e20d_return_output;
     VAR_printf_uxn_opcodes_h_l2730_c3_5f91_uxn_opcodes_h_l2730_c3_5f91_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2729_c1_cf07_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2754_c7_0dfe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;
     -- t8_MUX[uxn_opcodes_h_l2735_c7_652c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2735_c7_652c_cond <= VAR_t8_MUX_uxn_opcodes_h_l2735_c7_652c_cond;
     t8_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue;
     t8_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2735_c7_652c_return_output := t8_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2748_c7_e6b6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output;

     -- printf_uxn_opcodes_h_l2730_c3_5f91[uxn_opcodes_h_l2730_c3_5f91] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2730_c3_5f91_uxn_opcodes_h_l2730_c3_5f91_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2730_c3_5f91_uxn_opcodes_h_l2730_c3_5f91_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2744_c7_3775] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2744_c7_3775] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2748_c7_e6b6] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2735_c7_652c] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2744_c7_3775] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_return_output := result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;

     -- MUX[uxn_opcodes_h_l2742_c32_63d3] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2742_c32_63d3_cond <= VAR_MUX_uxn_opcodes_h_l2742_c32_63d3_cond;
     MUX_uxn_opcodes_h_l2742_c32_63d3_iftrue <= VAR_MUX_uxn_opcodes_h_l2742_c32_63d3_iftrue;
     MUX_uxn_opcodes_h_l2742_c32_63d3_iffalse <= VAR_MUX_uxn_opcodes_h_l2742_c32_63d3_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2742_c32_63d3_return_output := MUX_uxn_opcodes_h_l2742_c32_63d3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2748_c7_e6b6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue := VAR_MUX_uxn_opcodes_h_l2742_c32_63d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2748_c7_e6b6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;
     -- result_stack_value_MUX[uxn_opcodes_h_l2738_c7_1f6e] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output := result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2744_c7_3775] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;

     -- t8_MUX[uxn_opcodes_h_l2729_c2_ea1b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond <= VAR_t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond;
     t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue;
     t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output := t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2738_c7_1f6e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2738_c7_1f6e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2744_c7_3775] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2738_c7_1f6e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2744_c7_3775] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2729_c2_ea1b] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2744_c7_3775_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2735_c7_652c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2735_c7_652c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2738_c7_1f6e] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2738_c7_1f6e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2735_c7_652c] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_return_output := result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2735_c7_652c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2738_c7_1f6e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_1f6e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2729_c2_ea1b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2735_c7_652c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2729_c2_ea1b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2735_c7_652c] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2729_c2_ea1b] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output := result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2729_c2_ea1b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2735_c7_652c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2735_c7_652c_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2729_c2_ea1b] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2729_c2_ea1b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2729_c2_ea1b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_f6cd_uxn_opcodes_h_l2760_l2725_DUPLICATE_924a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f6cd_uxn_opcodes_h_l2760_l2725_DUPLICATE_924a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_f6cd(
     result,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2729_c2_ea1b_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f6cd_uxn_opcodes_h_l2760_l2725_DUPLICATE_924a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f6cd_uxn_opcodes_h_l2760_l2725_DUPLICATE_924a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
