-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity dup_0CLK_66ba3dc0 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_66ba3dc0;
architecture arch of dup_0CLK_66ba3dc0 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l3033_c6_80c1]
signal BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l3033_c1_e489]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l3033_c2_75cd]
signal t8_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3033_c2_75cd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3033_c2_75cd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3033_c2_75cd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l3033_c2_75cd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3033_c2_75cd]
signal result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3033_c2_75cd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l3034_c3_133c[uxn_opcodes_h_l3034_c3_133c]
signal printf_uxn_opcodes_h_l3034_c3_133c_uxn_opcodes_h_l3034_c3_133c_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3038_c11_5595]
signal BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l3038_c7_1560]
signal t8_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3038_c7_1560]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3038_c7_1560]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3038_c7_1560]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l3038_c7_1560]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3038_c7_1560]
signal result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3038_c7_1560]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3041_c11_df92]
signal BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l3041_c7_a6ee]
signal t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3041_c7_a6ee]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3041_c7_a6ee]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3041_c7_a6ee]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l3041_c7_a6ee]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3041_c7_a6ee]
signal result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3041_c7_a6ee]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l3044_c32_733a]
signal BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l3044_c32_89a0]
signal BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l3044_c32_8f3d]
signal MUX_uxn_opcodes_h_l3044_c32_8f3d_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l3044_c32_8f3d_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l3044_c32_8f3d_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l3044_c32_8f3d_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3046_c11_b7d1]
signal BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3046_c7_1dd9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3046_c7_1dd9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3046_c7_1dd9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3046_c7_1dd9]
signal result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3046_c7_1dd9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3052_c11_91f9]
signal BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3052_c7_9f51]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3052_c7_9f51]
signal result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3052_c7_9f51]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3052_c7_9f51]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3056_c11_06a5]
signal BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3056_c7_c68f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3056_c7_c68f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_09c5( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.stack_value := ref_toks_5;
      base.is_opc_done := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1
BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_left,
BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_right,
BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_return_output);

-- t8_MUX_uxn_opcodes_h_l3033_c2_75cd
t8_MUX_uxn_opcodes_h_l3033_c2_75cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l3033_c2_75cd_cond,
t8_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue,
t8_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse,
t8_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd
result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd
result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd
result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd
result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_cond,
result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd
result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output);

-- printf_uxn_opcodes_h_l3034_c3_133c_uxn_opcodes_h_l3034_c3_133c
printf_uxn_opcodes_h_l3034_c3_133c_uxn_opcodes_h_l3034_c3_133c : entity work.printf_uxn_opcodes_h_l3034_c3_133c_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l3034_c3_133c_uxn_opcodes_h_l3034_c3_133c_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595
BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_left,
BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_right,
BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_return_output);

-- t8_MUX_uxn_opcodes_h_l3038_c7_1560
t8_MUX_uxn_opcodes_h_l3038_c7_1560 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l3038_c7_1560_cond,
t8_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue,
t8_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse,
t8_MUX_uxn_opcodes_h_l3038_c7_1560_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560
result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560
result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560
result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560
result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_cond,
result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560
result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92
BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_left,
BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_right,
BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_return_output);

-- t8_MUX_uxn_opcodes_h_l3041_c7_a6ee
t8_MUX_uxn_opcodes_h_l3041_c7_a6ee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond,
t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue,
t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse,
t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee
result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee
result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee
result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee
result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond,
result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee
result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a
BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_left,
BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_right,
BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0
BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_left,
BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_right,
BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_return_output);

-- MUX_uxn_opcodes_h_l3044_c32_8f3d
MUX_uxn_opcodes_h_l3044_c32_8f3d : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l3044_c32_8f3d_cond,
MUX_uxn_opcodes_h_l3044_c32_8f3d_iftrue,
MUX_uxn_opcodes_h_l3044_c32_8f3d_iffalse,
MUX_uxn_opcodes_h_l3044_c32_8f3d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1
BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_left,
BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_right,
BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9
result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9
result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9
result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond,
result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9
result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9
BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_left,
BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_right,
BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51
result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_cond,
result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5
BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_left,
BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_right,
BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f
result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f
result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_return_output,
 t8_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_return_output,
 t8_MUX_uxn_opcodes_h_l3038_c7_1560_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_return_output,
 t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output,
 BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_return_output,
 BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_return_output,
 MUX_uxn_opcodes_h_l3044_c32_8f3d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3035_c3_cb46 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l3034_c3_133c_uxn_opcodes_h_l3034_c3_133c_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3039_c3_fd99 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3044_c32_8f3d_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3044_c32_8f3d_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3044_c32_8f3d_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3044_c32_8f3d_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3049_c3_4f26 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3053_c3_f9f8 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3033_l3056_l3052_l3041_l3038_DUPLICATE_373b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3033_l3046_l3038_DUPLICATE_35cf_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3041_l3033_l3038_DUPLICATE_d246_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3041_l3033_l3038_l3052_DUPLICATE_5075_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3056_l3052_l3046_l3041_l3038_DUPLICATE_8ab5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3041_l3052_DUPLICATE_de74_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_09c5_uxn_opcodes_h_l3061_l3029_DUPLICATE_4563_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3053_c3_f9f8 := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3053_c3_f9f8;
     VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3049_c3_4f26 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3049_c3_4f26;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_right := to_unsigned(5, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3039_c3_fd99 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3039_c3_fd99;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_right := to_unsigned(2, 2);
     VAR_MUX_uxn_opcodes_h_l3044_c32_8f3d_iffalse := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_right := to_unsigned(128, 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_iffalse := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l3044_c32_8f3d_iftrue := signed(std_logic_vector(resize(to_unsigned(2, 2), 8)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3035_c3_cb46 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3035_c3_cb46;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue := t8;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l3046_c11_b7d1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_left;
     BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_return_output := BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l3044_c32_733a] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_left;
     BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_return_output := BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3056_l3052_l3046_l3041_l3038_DUPLICATE_8ab5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3056_l3052_l3046_l3041_l3038_DUPLICATE_8ab5_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3033_l3046_l3038_DUPLICATE_35cf LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3033_l3046_l3038_DUPLICATE_35cf_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l3038_c11_5595] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_left;
     BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_return_output := BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l3033_c6_80c1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_left;
     BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output := BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l3052_c11_91f9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_left;
     BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_return_output := BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3041_l3033_l3038_l3052_DUPLICATE_5075 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3041_l3033_l3038_l3052_DUPLICATE_5075_return_output := result.stack_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l3056_c11_06a5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_left;
     BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_return_output := BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3041_l3052_DUPLICATE_de74 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3041_l3052_DUPLICATE_de74_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l3041_c11_df92] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_left;
     BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_return_output := BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3033_l3056_l3052_l3041_l3038_DUPLICATE_373b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3033_l3056_l3052_l3041_l3038_DUPLICATE_373b_return_output := result.is_stack_write;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3041_l3033_l3038_DUPLICATE_d246 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3041_l3033_l3038_DUPLICATE_d246_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_left := VAR_BIN_OP_AND_uxn_opcodes_h_l3044_c32_733a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3033_c6_80c1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3038_c7_1560_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3038_c11_5595_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3041_c11_df92_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3046_c11_b7d1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3052_c11_91f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3056_c11_06a5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3041_l3033_l3038_DUPLICATE_d246_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3041_l3033_l3038_DUPLICATE_d246_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3041_l3033_l3038_DUPLICATE_d246_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3056_l3052_l3046_l3041_l3038_DUPLICATE_8ab5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3056_l3052_l3046_l3041_l3038_DUPLICATE_8ab5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3056_l3052_l3046_l3041_l3038_DUPLICATE_8ab5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3056_l3052_l3046_l3041_l3038_DUPLICATE_8ab5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3056_l3052_l3046_l3041_l3038_DUPLICATE_8ab5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3033_l3046_l3038_DUPLICATE_35cf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3033_l3046_l3038_DUPLICATE_35cf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3033_l3046_l3038_DUPLICATE_35cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3033_l3056_l3052_l3041_l3038_DUPLICATE_373b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3033_l3056_l3052_l3041_l3038_DUPLICATE_373b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3033_l3056_l3052_l3041_l3038_DUPLICATE_373b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3033_l3056_l3052_l3041_l3038_DUPLICATE_373b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3033_l3056_l3052_l3041_l3038_DUPLICATE_373b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3041_l3052_DUPLICATE_de74_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3041_l3052_DUPLICATE_de74_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3041_l3033_l3038_l3052_DUPLICATE_5075_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3041_l3033_l3038_l3052_DUPLICATE_5075_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3041_l3033_l3038_l3052_DUPLICATE_5075_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3041_l3033_l3038_l3052_DUPLICATE_5075_return_output;
     -- t8_MUX[uxn_opcodes_h_l3041_c7_a6ee] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond <= VAR_t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond;
     t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue;
     t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output := t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3056_c7_c68f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3056_c7_c68f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3052_c7_9f51] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output := result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3046_c7_1dd9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l3044_c32_89a0] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_left;
     BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_return_output := BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3052_c7_9f51] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l3033_c1_e489] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l3044_c32_8f3d_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l3044_c32_89a0_return_output;
     VAR_printf_uxn_opcodes_h_l3034_c3_133c_uxn_opcodes_h_l3034_c3_133c_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3033_c1_e489_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3056_c7_c68f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse := VAR_t8_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;
     -- t8_MUX[uxn_opcodes_h_l3038_c7_1560] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l3038_c7_1560_cond <= VAR_t8_MUX_uxn_opcodes_h_l3038_c7_1560_cond;
     t8_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue;
     t8_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l3038_c7_1560_return_output := t8_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3052_c7_9f51] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3046_c7_1dd9] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output := result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3046_c7_1dd9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3041_c7_a6ee] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;

     -- printf_uxn_opcodes_h_l3034_c3_133c[uxn_opcodes_h_l3034_c3_133c] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l3034_c3_133c_uxn_opcodes_h_l3034_c3_133c_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l3034_c3_133c_uxn_opcodes_h_l3034_c3_133c_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- MUX[uxn_opcodes_h_l3044_c32_8f3d] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l3044_c32_8f3d_cond <= VAR_MUX_uxn_opcodes_h_l3044_c32_8f3d_cond;
     MUX_uxn_opcodes_h_l3044_c32_8f3d_iftrue <= VAR_MUX_uxn_opcodes_h_l3044_c32_8f3d_iftrue;
     MUX_uxn_opcodes_h_l3044_c32_8f3d_iffalse <= VAR_MUX_uxn_opcodes_h_l3044_c32_8f3d_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l3044_c32_8f3d_return_output := MUX_uxn_opcodes_h_l3044_c32_8f3d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3052_c7_9f51] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue := VAR_MUX_uxn_opcodes_h_l3044_c32_8f3d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3052_c7_9f51_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse := VAR_t8_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;
     -- t8_MUX[uxn_opcodes_h_l3033_c2_75cd] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l3033_c2_75cd_cond <= VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75cd_cond;
     t8_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue;
     t8_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output := t8_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3041_c7_a6ee] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3041_c7_a6ee] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output := result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l3041_c7_a6ee] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3046_c7_1dd9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3038_c7_1560] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3046_c7_1dd9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3046_c7_1dd9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output;
     -- result_stack_value_MUX[uxn_opcodes_h_l3038_c7_1560] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_return_output := result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3041_c7_a6ee] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3041_c7_a6ee] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3038_c7_1560] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l3038_c7_1560] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3033_c2_75cd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3041_c7_a6ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l3038_c7_1560] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3033_c2_75cd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l3033_c2_75cd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3038_c7_1560] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3033_c2_75cd] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output := result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3038_c7_1560_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l3033_c2_75cd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3033_c2_75cd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_09c5_uxn_opcodes_h_l3061_l3029_DUPLICATE_4563 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_09c5_uxn_opcodes_h_l3061_l3029_DUPLICATE_4563_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_09c5(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3033_c2_75cd_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_09c5_uxn_opcodes_h_l3061_l3029_DUPLICATE_4563_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_09c5_uxn_opcodes_h_l3061_l3029_DUPLICATE_4563_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
