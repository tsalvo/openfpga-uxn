-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity sub1_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub1_0CLK_64d180f1;
architecture arch of sub1_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2461_c6_d6a5]
signal BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2461_c2_9edf]
signal t8_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2461_c2_9edf]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2461_c2_9edf]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2461_c2_9edf]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2461_c2_9edf]
signal result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2461_c2_9edf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2461_c2_9edf]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2461_c2_9edf]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2461_c2_9edf]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2461_c2_9edf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2461_c2_9edf]
signal n8_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2474_c11_73c3]
signal BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2474_c7_ea0f]
signal t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2474_c7_ea0f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2474_c7_ea0f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2474_c7_ea0f]
signal result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2474_c7_ea0f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2474_c7_ea0f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2474_c7_ea0f]
signal n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2477_c11_f671]
signal BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2477_c7_4076]
signal t8_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2477_c7_4076]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2477_c7_4076]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2477_c7_4076]
signal result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2477_c7_4076]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2477_c7_4076]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2477_c7_4076]
signal n8_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2480_c11_9156]
signal BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2480_c7_9450]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2480_c7_9450]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2480_c7_9450]
signal result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2480_c7_9450]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2480_c7_9450]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2480_c7_9450]
signal n8_MUX_uxn_opcodes_h_l2480_c7_9450_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2480_c7_9450_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2482_c30_1a2b]
signal sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_return_output : signed(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2485_c21_5d97]
signal BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_71f0( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_index_flipped := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5
BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_left,
BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_right,
BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output);

-- t8_MUX_uxn_opcodes_h_l2461_c2_9edf
t8_MUX_uxn_opcodes_h_l2461_c2_9edf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2461_c2_9edf_cond,
t8_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue,
t8_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse,
t8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_cond,
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output);

-- n8_MUX_uxn_opcodes_h_l2461_c2_9edf
n8_MUX_uxn_opcodes_h_l2461_c2_9edf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2461_c2_9edf_cond,
n8_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue,
n8_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse,
n8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3
BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_left,
BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_right,
BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_return_output);

-- t8_MUX_uxn_opcodes_h_l2474_c7_ea0f
t8_MUX_uxn_opcodes_h_l2474_c7_ea0f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond,
t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue,
t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse,
t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output);

-- n8_MUX_uxn_opcodes_h_l2474_c7_ea0f
n8_MUX_uxn_opcodes_h_l2474_c7_ea0f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond,
n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue,
n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse,
n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671
BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_left,
BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_right,
BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_return_output);

-- t8_MUX_uxn_opcodes_h_l2477_c7_4076
t8_MUX_uxn_opcodes_h_l2477_c7_4076 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2477_c7_4076_cond,
t8_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue,
t8_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse,
t8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_cond,
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_return_output);

-- n8_MUX_uxn_opcodes_h_l2477_c7_4076
n8_MUX_uxn_opcodes_h_l2477_c7_4076 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2477_c7_4076_cond,
n8_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue,
n8_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse,
n8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156
BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_left,
BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_right,
BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_cond,
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_return_output);

-- n8_MUX_uxn_opcodes_h_l2480_c7_9450
n8_MUX_uxn_opcodes_h_l2480_c7_9450 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2480_c7_9450_cond,
n8_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue,
n8_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse,
n8_MUX_uxn_opcodes_h_l2480_c7_9450_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b
sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_ins,
sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_x,
sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_y,
sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97
BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_left,
BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_right,
BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output,
 t8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
 n8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_return_output,
 t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output,
 n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_return_output,
 t8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_return_output,
 n8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_return_output,
 n8_MUX_uxn_opcodes_h_l2480_c7_9450_return_output,
 sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2466_c3_f9c8 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2471_c3_507a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2461_c2_9edf_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2475_c3_69ac : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2480_c7_9450_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2477_c7_4076_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2484_c3_ff00 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2480_c7_9450_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2461_l2480_l2474_l2477_DUPLICATE_fb5e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_07c4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_01e8_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_04a9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2480_l2477_DUPLICATE_085e_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2489_l2457_DUPLICATE_650d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2466_c3_f9c8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2466_c3_f9c8;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2475_c3_69ac := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2475_c3_69ac;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2484_c3_ff00 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2484_c3_ff00;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2471_c3_507a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2471_c3_507a;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2480_c11_9156] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_left;
     BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_return_output := BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2461_c2_9edf_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2474_c11_73c3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_left;
     BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_return_output := BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2461_c2_9edf_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2480_l2477_DUPLICATE_085e LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2480_l2477_DUPLICATE_085e_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2461_c2_9edf_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_01e8 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_01e8_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_04a9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_04a9_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2461_c6_d6a5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2482_c30_1a2b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_ins;
     sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_x;
     sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_return_output := sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_return_output;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2485_c21_5d97] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2461_c2_9edf_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2461_l2480_l2474_l2477_DUPLICATE_fb5e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2461_l2480_l2474_l2477_DUPLICATE_fb5e_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_07c4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_07c4_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2477_c11_f671] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_left;
     BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_return_output := BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2461_c2_9edf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2461_c2_9edf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2461_c6_d6a5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2474_c11_73c3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2477_c7_4076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2477_c7_4076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2477_c11_f671_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2480_c7_9450_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2480_c11_9156_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2485_c21_5d97_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_01e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_01e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_01e8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_04a9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_04a9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_04a9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_07c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_07c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2480_l2474_l2477_DUPLICATE_07c4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2480_l2477_DUPLICATE_085e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2480_l2477_DUPLICATE_085e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2461_l2480_l2474_l2477_DUPLICATE_fb5e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2461_l2480_l2474_l2477_DUPLICATE_fb5e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2461_l2480_l2474_l2477_DUPLICATE_fb5e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2461_l2480_l2474_l2477_DUPLICATE_fb5e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2461_c2_9edf_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2461_c2_9edf_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2461_c2_9edf_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2461_c2_9edf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2482_c30_1a2b_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2480_c7_9450] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2480_c7_9450] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2480_c7_9450] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2480_c7_9450] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output;

     -- n8_MUX[uxn_opcodes_h_l2480_c7_9450] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2480_c7_9450_cond <= VAR_n8_MUX_uxn_opcodes_h_l2480_c7_9450_cond;
     n8_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue;
     n8_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2480_c7_9450_return_output := n8_MUX_uxn_opcodes_h_l2480_c7_9450_return_output;

     -- t8_MUX[uxn_opcodes_h_l2477_c7_4076] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2477_c7_4076_cond <= VAR_t8_MUX_uxn_opcodes_h_l2477_c7_4076_cond;
     t8_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue;
     t8_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output := t8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2480_c7_9450] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_return_output := result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2480_c7_9450_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2480_c7_9450_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2480_c7_9450_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2480_c7_9450_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2480_c7_9450_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2480_c7_9450_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2477_c7_4076] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2477_c7_4076] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_return_output := result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;

     -- t8_MUX[uxn_opcodes_h_l2474_c7_ea0f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond;
     t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue;
     t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output := t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2477_c7_4076] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;

     -- n8_MUX[uxn_opcodes_h_l2477_c7_4076] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2477_c7_4076_cond <= VAR_n8_MUX_uxn_opcodes_h_l2477_c7_4076_cond;
     n8_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue;
     n8_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output := n8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2477_c7_4076] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2477_c7_4076] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2477_c7_4076_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;
     -- t8_MUX[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2461_c2_9edf_cond <= VAR_t8_MUX_uxn_opcodes_h_l2461_c2_9edf_cond;
     t8_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue;
     t8_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output := t8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output;

     -- n8_MUX[uxn_opcodes_h_l2474_c7_ea0f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond;
     n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue;
     n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output := n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2474_c7_ea0f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2474_c7_ea0f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2474_c7_ea0f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2474_c7_ea0f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2474_c7_ea0f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2474_c7_ea0f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output;

     -- n8_MUX[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2461_c2_9edf_cond <= VAR_n8_MUX_uxn_opcodes_h_l2461_c2_9edf_cond;
     n8_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue;
     n8_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output := n8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2461_c2_9edf] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output := result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2489_l2457_DUPLICATE_650d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2489_l2457_DUPLICATE_650d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_71f0(
     result,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2461_c2_9edf_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2489_l2457_DUPLICATE_650d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2489_l2457_DUPLICATE_650d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
