-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 57
entity nip2_0CLK_4dee2d7a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_4dee2d7a;
architecture arch of nip2_0CLK_4dee2d7a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2310_c6_36bd]
signal BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2310_c2_f8b7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2310_c2_f8b7]
signal result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2310_c2_f8b7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2310_c2_f8b7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2310_c2_f8b7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2310_c2_f8b7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2310_c2_f8b7]
signal t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2315_c11_9f8d]
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2315_c7_a412]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2315_c7_a412]
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2315_c7_a412]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2315_c7_a412]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2315_c7_a412]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2315_c7_a412]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2315_c7_a412]
signal t16_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2318_c11_73f2]
signal BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2318_c7_4b60]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2318_c7_4b60]
signal result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2318_c7_4b60]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2318_c7_4b60]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2318_c7_4b60]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2318_c7_4b60]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2318_c7_4b60]
signal t16_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2320_c3_bff5]
signal CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2323_c11_00cf]
signal BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2323_c7_89c3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2323_c7_89c3]
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2323_c7_89c3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2323_c7_89c3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2323_c7_89c3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2323_c7_89c3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2323_c7_89c3]
signal t16_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2326_c11_2349]
signal BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2326_c7_90c8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2326_c7_90c8]
signal result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2326_c7_90c8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2326_c7_90c8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2326_c7_90c8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2326_c7_90c8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2326_c7_90c8]
signal t16_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2327_c3_0666]
signal BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2329_c30_e63c]
signal sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2334_c11_09e8]
signal BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2334_c7_effe]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2334_c7_effe]
signal result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2334_c7_effe]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2334_c7_effe]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2334_c7_effe]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_return_output : unsigned(0 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l2337_c31_aba0]
signal CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2339_c11_e01f]
signal BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2339_c7_98a9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2339_c7_98a9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_3345( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd
BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_left,
BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_right,
BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7
result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond,
result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7
result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7
result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7
result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7
result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output);

-- t16_MUX_uxn_opcodes_h_l2310_c2_f8b7
t16_MUX_uxn_opcodes_h_l2310_c2_f8b7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond,
t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue,
t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse,
t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_left,
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_right,
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_cond,
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412
result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output);

-- t16_MUX_uxn_opcodes_h_l2315_c7_a412
t16_MUX_uxn_opcodes_h_l2315_c7_a412 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2315_c7_a412_cond,
t16_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue,
t16_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse,
t16_MUX_uxn_opcodes_h_l2315_c7_a412_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2
BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_left,
BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_right,
BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60
result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_cond,
result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60
result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60
result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60
result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60
result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output);

-- t16_MUX_uxn_opcodes_h_l2318_c7_4b60
t16_MUX_uxn_opcodes_h_l2318_c7_4b60 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2318_c7_4b60_cond,
t16_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue,
t16_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse,
t16_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5
CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5_x,
CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_left,
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_right,
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3
result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3
result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output);

-- t16_MUX_uxn_opcodes_h_l2323_c7_89c3
t16_MUX_uxn_opcodes_h_l2323_c7_89c3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2323_c7_89c3_cond,
t16_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue,
t16_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse,
t16_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349
BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_left,
BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_right,
BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8
result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8
result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8
result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8
result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output);

-- t16_MUX_uxn_opcodes_h_l2326_c7_90c8
t16_MUX_uxn_opcodes_h_l2326_c7_90c8 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2326_c7_90c8_cond,
t16_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue,
t16_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse,
t16_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666
BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_left,
BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_right,
BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c
sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_ins,
sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_x,
sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_y,
sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8
BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_left,
BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_right,
BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe
result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_cond,
result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe
result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe
result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe
result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_return_output);

-- CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0
CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0_x,
CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f
BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_left,
BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_right,
BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9
result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output,
 t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output,
 t16_MUX_uxn_opcodes_h_l2315_c7_a412_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output,
 t16_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output,
 CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output,
 t16_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output,
 t16_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_return_output,
 sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_return_output,
 CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2312_c3_07fd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_a412_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2316_c3_134a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_a412_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2321_c3_1408 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2318_c7_4b60_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2324_c3_bf44 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2323_c7_89c3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2331_c3_9079 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2326_c7_90c8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_return_output : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2332_c21_1cde_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2336_c3_425e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2334_c7_effe_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2337_c21_93aa_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b09c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2339_l2310_DUPLICATE_89d9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2326_l2323_l2318_l2315_l2310_DUPLICATE_1336_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b059_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2334_l2326_l2323_l2318_l2315_l2339_DUPLICATE_a930_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2319_l2327_DUPLICATE_c5e3_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2306_l2344_DUPLICATE_7c0c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_y := resize(to_signed(-2, 3), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2316_c3_134a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2316_c3_134a;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2336_c3_425e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2336_c3_425e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2321_c3_1408 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2321_c3_1408;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_right := to_unsigned(6, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2331_c3_9079 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2331_c3_9079;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2312_c3_07fd := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2312_c3_07fd;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2324_c3_bf44 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2324_c3_bf44;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_left := t16;
     VAR_CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0_x := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse := t16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b059 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b059_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2326_c11_2349] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_left;
     BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_return_output := BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2329_c30_e63c] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_ins;
     sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_x;
     sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_return_output := sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2315_c11_9f8d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2339_c11_e01f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2334_c7_effe] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2334_c7_effe_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2326_l2323_l2318_l2315_l2310_DUPLICATE_1336 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2326_l2323_l2318_l2315_l2310_DUPLICATE_1336_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2323_c11_00cf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_left;
     BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_return_output := BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_return_output;

     -- CONST_SR_8[uxn_opcodes_h_l2337_c31_aba0] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0_x <= VAR_CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0_return_output := CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2334_c11_09e8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2334_l2326_l2323_l2318_l2315_l2339_DUPLICATE_a930 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2334_l2326_l2323_l2318_l2315_l2339_DUPLICATE_a930_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2310_c6_36bd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2319_l2327_DUPLICATE_c5e3 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2319_l2327_DUPLICATE_c5e3_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l2318_c11_73f2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b09c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b09c_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2339_l2310_DUPLICATE_89d9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2339_l2310_DUPLICATE_89d9_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2310_c6_36bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_a412_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_9f8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2318_c7_4b60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2318_c11_73f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2323_c7_89c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_00cf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2326_c7_90c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2326_c11_2349_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2334_c11_09e8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_e01f_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2319_l2327_DUPLICATE_c5e3_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2319_l2327_DUPLICATE_c5e3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2326_l2323_l2318_l2315_l2310_DUPLICATE_1336_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2326_l2323_l2318_l2315_l2310_DUPLICATE_1336_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2326_l2323_l2318_l2315_l2310_DUPLICATE_1336_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2326_l2323_l2318_l2315_l2310_DUPLICATE_1336_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2326_l2323_l2318_l2315_l2310_DUPLICATE_1336_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2334_l2326_l2323_l2318_l2315_l2339_DUPLICATE_a930_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2334_l2326_l2323_l2318_l2315_l2339_DUPLICATE_a930_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2334_l2326_l2323_l2318_l2315_l2339_DUPLICATE_a930_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2334_l2326_l2323_l2318_l2315_l2339_DUPLICATE_a930_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2334_l2326_l2323_l2318_l2315_l2339_DUPLICATE_a930_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2334_l2326_l2323_l2318_l2315_l2339_DUPLICATE_a930_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b059_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b059_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b059_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b059_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b059_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2339_l2310_DUPLICATE_89d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2339_l2310_DUPLICATE_89d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2339_l2310_DUPLICATE_89d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2339_l2310_DUPLICATE_89d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2339_l2310_DUPLICATE_89d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2339_l2310_DUPLICATE_89d9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b09c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b09c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b09c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b09c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2334_l2323_l2318_l2315_l2310_DUPLICATE_b09c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2334_c7_effe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2329_c30_e63c_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2326_c7_90c8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2334_c7_effe] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2339_c7_98a9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2339_c7_98a9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2337_c21_93aa] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2337_c21_93aa_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l2337_c31_aba0_return_output);

     -- CONST_SL_8[uxn_opcodes_h_l2320_c3_bff5] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5_return_output := CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2327_c3_0666] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_left;
     BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_return_output := BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2334_c7_effe] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2337_c21_93aa_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2320_c3_bff5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2334_c7_effe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2339_c7_98a9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2334_c7_effe_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2326_c7_90c8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2332_c21_1cde] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2332_c21_1cde_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_BIN_OP_OR_uxn_opcodes_h_l2327_c3_0666_return_output);

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2334_c7_effe] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2334_c7_effe] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_return_output := result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2334_c7_effe] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_return_output;

     -- t16_MUX[uxn_opcodes_h_l2326_c7_90c8] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2326_c7_90c8_cond <= VAR_t16_MUX_uxn_opcodes_h_l2326_c7_90c8_cond;
     t16_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue;
     t16_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output := t16_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2323_c7_89c3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2326_c7_90c8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2332_c21_1cde_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2334_c7_effe_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2334_c7_effe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2334_c7_effe_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2326_c7_90c8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2323_c7_89c3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;

     -- t16_MUX[uxn_opcodes_h_l2323_c7_89c3] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2323_c7_89c3_cond <= VAR_t16_MUX_uxn_opcodes_h_l2323_c7_89c3_cond;
     t16_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue;
     t16_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output := t16_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2318_c7_4b60] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2326_c7_90c8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2326_c7_90c8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2323_c7_89c3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2326_c7_90c8_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2323_c7_89c3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2318_c7_4b60] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2318_c7_4b60] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2323_c7_89c3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2315_c7_a412] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2323_c7_89c3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;

     -- t16_MUX[uxn_opcodes_h_l2318_c7_4b60] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2318_c7_4b60_cond <= VAR_t16_MUX_uxn_opcodes_h_l2318_c7_4b60_cond;
     t16_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue;
     t16_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output := t16_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_89c3_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;
     -- t16_MUX[uxn_opcodes_h_l2315_c7_a412] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2315_c7_a412_cond <= VAR_t16_MUX_uxn_opcodes_h_l2315_c7_a412_cond;
     t16_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue;
     t16_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_a412_return_output := t16_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2310_c2_f8b7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2318_c7_4b60] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2315_c7_a412] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2318_c7_4b60] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2318_c7_4b60] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output := result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2315_c7_a412] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2318_c7_4b60_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2310_c2_f8b7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2310_c2_f8b7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output;

     -- t16_MUX[uxn_opcodes_h_l2310_c2_f8b7] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond <= VAR_t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond;
     t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue;
     t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output := t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2315_c7_a412] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_return_output := result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2315_c7_a412] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2315_c7_a412] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_a412_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2310_c2_f8b7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2310_c2_f8b7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2310_c2_f8b7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output := result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2306_l2344_DUPLICATE_7c0c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2306_l2344_DUPLICATE_7c0c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3345(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2310_c2_f8b7_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2306_l2344_DUPLICATE_7c0c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2306_l2344_DUPLICATE_7c0c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
