-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sft_0CLK_8d2aa467 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sft_0CLK_8d2aa467;
architecture arch of sft_0CLK_8d2aa467 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2213_c6_1efb]
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2213_c2_ec4e]
signal n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2213_c2_ec4e]
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2213_c2_ec4e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2213_c2_ec4e]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2213_c2_ec4e]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2213_c2_ec4e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2213_c2_ec4e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2213_c2_ec4e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2213_c2_ec4e]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2213_c2_ec4e]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2213_c2_ec4e]
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2213_c2_ec4e]
signal t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2226_c11_ee16]
signal BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2226_c7_81ff]
signal n8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2226_c7_81ff]
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2226_c7_81ff]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2226_c7_81ff]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2226_c7_81ff]
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2226_c7_81ff]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2226_c7_81ff]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2226_c7_81ff]
signal t8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2229_c11_6b10]
signal BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2229_c7_f98f]
signal n8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2229_c7_f98f]
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2229_c7_f98f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2229_c7_f98f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2229_c7_f98f]
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2229_c7_f98f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2229_c7_f98f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2229_c7_f98f]
signal t8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2231_c30_33a3]
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2233_c11_ffdd]
signal BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2233_c7_8eb2]
signal n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2233_c7_8eb2]
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2233_c7_8eb2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2233_c7_8eb2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2233_c7_8eb2]
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2233_c7_8eb2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2233_c7_8eb2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2236_c18_3c39]
signal BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_return_output : unsigned(7 downto 0);

-- BIN_OP_SR[uxn_opcodes_h_l2236_c11_87b2]
signal BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_left : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_right : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_return_output : unsigned(7 downto 0);

-- CONST_SR_4[uxn_opcodes_h_l2236_c34_6962]
signal CONST_SR_4_uxn_opcodes_h_l2236_c34_6962_x : unsigned(7 downto 0);
signal CONST_SR_4_uxn_opcodes_h_l2236_c34_6962_return_output : unsigned(7 downto 0);

-- BIN_OP_SL[uxn_opcodes_h_l2236_c11_6d0f]
signal BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_left : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_right : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8b52( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_left,
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_right,
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output);

-- n8_MUX_uxn_opcodes_h_l2213_c2_ec4e
n8_MUX_uxn_opcodes_h_l2213_c2_ec4e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond,
n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue,
n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse,
n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e
tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond,
tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue,
tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse,
tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output);

-- t8_MUX_uxn_opcodes_h_l2213_c2_ec4e
t8_MUX_uxn_opcodes_h_l2213_c2_ec4e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond,
t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue,
t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse,
t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_left,
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_right,
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output);

-- n8_MUX_uxn_opcodes_h_l2226_c7_81ff
n8_MUX_uxn_opcodes_h_l2226_c7_81ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond,
n8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue,
n8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse,
n8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff
tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond,
tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue,
tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse,
tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_cond,
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output);

-- t8_MUX_uxn_opcodes_h_l2226_c7_81ff
t8_MUX_uxn_opcodes_h_l2226_c7_81ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond,
t8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue,
t8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse,
t8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_left,
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_right,
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output);

-- n8_MUX_uxn_opcodes_h_l2229_c7_f98f
n8_MUX_uxn_opcodes_h_l2229_c7_f98f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond,
n8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue,
n8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse,
n8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f
tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond,
tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue,
tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse,
tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output);

-- t8_MUX_uxn_opcodes_h_l2229_c7_f98f
t8_MUX_uxn_opcodes_h_l2229_c7_f98f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond,
t8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue,
t8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse,
t8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3
sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_ins,
sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_x,
sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_y,
sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_left,
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_right,
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_return_output);

-- n8_MUX_uxn_opcodes_h_l2233_c7_8eb2
n8_MUX_uxn_opcodes_h_l2233_c7_8eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond,
n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue,
n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse,
n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2
tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond,
tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue,
tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse,
tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39
BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_left,
BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_right,
BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_return_output);

-- BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2
BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2 : entity work.BIN_OP_SR_uint8_t_uint8_t_0CLK_41db8d51 port map (
BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_left,
BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_right,
BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_return_output);

-- CONST_SR_4_uxn_opcodes_h_l2236_c34_6962
CONST_SR_4_uxn_opcodes_h_l2236_c34_6962 : entity work.CONST_SR_4_uint8_t_0CLK_de264c78 port map (
CONST_SR_4_uxn_opcodes_h_l2236_c34_6962_x,
CONST_SR_4_uxn_opcodes_h_l2236_c34_6962_return_output);

-- BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f
BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f : entity work.BIN_OP_SL_uint8_t_uint8_t_0CLK_ad8922d4 port map (
BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_left,
BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_right,
BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output,
 n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
 tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
 t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output,
 n8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output,
 tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output,
 t8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output,
 n8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output,
 tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output,
 t8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output,
 sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_return_output,
 n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output,
 tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_return_output,
 BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_return_output,
 CONST_SR_4_uxn_opcodes_h_l2236_c34_6962_return_output,
 BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2218_c3_ec7d : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_ba79 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2227_c3_2d84 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_be4f : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2238_c3_5b09 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_left : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_6962_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_right : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_6962_x : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_1e2b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2226_l2233_DUPLICATE_dd1d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_b6d9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_e36d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_c84d_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2243_l2209_DUPLICATE_b250_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2218_c3_ec7d := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2218_c3_ec7d;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_right := to_unsigned(15, 8);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2227_c3_2d84 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2227_c3_2d84;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_be4f := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_be4f;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_ba79 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_ba79;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2238_c3_5b09 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2238_c3_5b09;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_left := VAR_phase;
     VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_left := t8;
     VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_6962_x := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2229_c11_6b10] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_left;
     BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output := BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2213_c6_1efb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_left;
     BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output := BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2233_c11_ffdd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2231_c30_33a3] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_ins;
     sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_x;
     sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_return_output := sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_b6d9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_b6d9_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_e36d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_e36d_return_output := result.is_opc_done;

     -- CONST_SR_4[uxn_opcodes_h_l2236_c34_6962] LATENCY=0
     -- Inputs
     CONST_SR_4_uxn_opcodes_h_l2236_c34_6962_x <= VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_6962_x;
     -- Outputs
     VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_6962_return_output := CONST_SR_4_uxn_opcodes_h_l2236_c34_6962_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2226_l2233_DUPLICATE_dd1d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2226_l2233_DUPLICATE_dd1d_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_1e2b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_1e2b_return_output := result.u8_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2213_c2_ec4e_return_output := result.is_ram_write;

     -- BIN_OP_AND[uxn_opcodes_h_l2236_c18_3c39] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_left;
     BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_return_output := BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2213_c2_ec4e_return_output := result.is_pc_updated;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2213_c2_ec4e_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_c84d LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_c84d_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2226_c11_ee16] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_left;
     BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output := BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2213_c2_ec4e_return_output := result.is_vram_write;

     -- Submodule level 1
     VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_right := VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_3c39_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1efb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_ee16_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_6b10_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_ffdd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2226_l2233_DUPLICATE_dd1d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2226_l2233_DUPLICATE_dd1d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_e36d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_e36d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_e36d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_b6d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_b6d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_b6d9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_c84d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_c84d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_1e2b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_1e2b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_1e2b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_1e2b_return_output;
     VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_right := VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_6962_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2213_c2_ec4e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2213_c2_ec4e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2213_c2_ec4e_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2213_c2_ec4e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_33a3_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2233_c7_8eb2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2233_c7_8eb2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;

     -- t8_MUX[uxn_opcodes_h_l2229_c7_f98f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond;
     t8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue;
     t8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output := t8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;

     -- n8_MUX[uxn_opcodes_h_l2233_c7_8eb2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond <= VAR_n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond;
     n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue;
     n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output := n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2233_c7_8eb2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;

     -- BIN_OP_SR[uxn_opcodes_h_l2236_c11_87b2] LATENCY=0
     -- Inputs
     BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_left <= VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_left;
     BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_right <= VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_right;
     -- Outputs
     VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_return_output := BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2233_c7_8eb2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;

     -- Submodule level 2
     VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_left := VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_87b2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2229_c7_f98f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;

     -- t8_MUX[uxn_opcodes_h_l2226_c7_81ff] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond <= VAR_t8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond;
     t8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue;
     t8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output := t8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2229_c7_f98f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2229_c7_f98f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;

     -- n8_MUX[uxn_opcodes_h_l2229_c7_f98f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond;
     n8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue;
     n8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output := n8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2229_c7_f98f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;

     -- BIN_OP_SL[uxn_opcodes_h_l2236_c11_6d0f] LATENCY=0
     -- Inputs
     BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_left <= VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_left;
     BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_right <= VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_right;
     -- Outputs
     VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_return_output := BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_6d0f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2226_c7_81ff] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2233_c7_8eb2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;

     -- t8_MUX[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond <= VAR_t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond;
     t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue;
     t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output := t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2226_c7_81ff] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond <= VAR_n8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond;
     n8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue;
     n8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output := n8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2226_c7_81ff] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2226_c7_81ff] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2233_c7_8eb2] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_cond;
     tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output := tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2226_c7_81ff] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_8eb2_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2229_c7_f98f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2229_c7_f98f] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_cond;
     tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output := tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond <= VAR_n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond;
     n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue;
     n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output := n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f98f_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2226_c7_81ff] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_cond;
     tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output := tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2226_c7_81ff] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output := result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_81ff_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2213_c2_ec4e] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_cond;
     tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output := tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;

     -- Submodule level 7
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2243_l2209_DUPLICATE_b250 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2243_l2209_DUPLICATE_b250_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8b52(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_ec4e_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2243_l2209_DUPLICATE_b250_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2243_l2209_DUPLICATE_b250_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
