-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 37
entity dup_0CLK_6be78140 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_6be78140;
architecture arch of dup_0CLK_6be78140 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2958_c6_0764]
signal BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2958_c1_f670]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2958_c2_de38]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2958_c2_de38]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2958_c2_de38]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2958_c2_de38]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2958_c2_de38]
signal result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2958_c2_de38]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2958_c2_de38]
signal t8_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2959_c3_147d[uxn_opcodes_h_l2959_c3_147d]
signal printf_uxn_opcodes_h_l2959_c3_147d_uxn_opcodes_h_l2959_c3_147d_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2963_c11_afb7]
signal BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2963_c7_6c80]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2963_c7_6c80]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2963_c7_6c80]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2963_c7_6c80]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2963_c7_6c80]
signal result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2963_c7_6c80]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2963_c7_6c80]
signal t8_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2966_c11_1428]
signal BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2966_c7_c3b2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2966_c7_c3b2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2966_c7_c3b2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2966_c7_c3b2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2966_c7_c3b2]
signal result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2966_c7_c3b2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2966_c7_c3b2]
signal t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2969_c30_056c]
signal sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2974_c11_5c5e]
signal BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2974_c7_a7ab]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2974_c7_a7ab]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2974_c7_a7ab]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2974_c7_a7ab]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2974_c7_a7ab]
signal result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2979_c11_a26a]
signal BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2979_c7_fd5f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2979_c7_fd5f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_641b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764
BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_left,
BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_right,
BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38
result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38
result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38
result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38
result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_cond,
result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38
result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output);

-- t8_MUX_uxn_opcodes_h_l2958_c2_de38
t8_MUX_uxn_opcodes_h_l2958_c2_de38 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2958_c2_de38_cond,
t8_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue,
t8_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse,
t8_MUX_uxn_opcodes_h_l2958_c2_de38_return_output);

-- printf_uxn_opcodes_h_l2959_c3_147d_uxn_opcodes_h_l2959_c3_147d
printf_uxn_opcodes_h_l2959_c3_147d_uxn_opcodes_h_l2959_c3_147d : entity work.printf_uxn_opcodes_h_l2959_c3_147d_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2959_c3_147d_uxn_opcodes_h_l2959_c3_147d_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7
BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_left,
BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_right,
BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80
result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80
result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80
result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80
result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_cond,
result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80
result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output);

-- t8_MUX_uxn_opcodes_h_l2963_c7_6c80
t8_MUX_uxn_opcodes_h_l2963_c7_6c80 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2963_c7_6c80_cond,
t8_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue,
t8_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse,
t8_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428
BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_left,
BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_right,
BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2
result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2
result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2
result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2
result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output);

-- t8_MUX_uxn_opcodes_h_l2966_c7_c3b2
t8_MUX_uxn_opcodes_h_l2966_c7_c3b2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond,
t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue,
t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse,
t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2969_c30_056c
sp_relative_shift_uxn_opcodes_h_l2969_c30_056c : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_ins,
sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_x,
sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_y,
sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e
BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_left,
BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_right,
BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab
result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab
result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab
result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab
result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond,
result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a
BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_left,
BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_right,
BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f
result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f
result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output,
 t8_MUX_uxn_opcodes_h_l2958_c2_de38_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output,
 t8_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output,
 t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output,
 sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2960_c3_274f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2958_c2_de38_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2958_c2_de38_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2959_c3_147d_uxn_opcodes_h_l2959_c3_147d_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2964_c3_567c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2963_c7_6c80_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2971_c3_05a4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2976_c3_b551 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2974_c7_a7ab_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2958_l2974_l2963_DUPLICATE_7517_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2958_l2974_l2963_l2979_DUPLICATE_b1c1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2958_l2974_l2963_DUPLICATE_e2fc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2958_l2963_l2966_DUPLICATE_4cb8_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2974_l2963_l2979_l2966_DUPLICATE_ba35_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2984_l2954_DUPLICATE_e679_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2964_c3_567c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2964_c3_567c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_right := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_iffalse := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2976_c3_b551 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2976_c3_b551;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2960_c3_274f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2960_c3_274f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2971_c3_05a4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2971_c3_05a4;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2966_c11_1428] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_left;
     BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_return_output := BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2958_l2963_l2966_DUPLICATE_4cb8 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2958_l2963_l2966_DUPLICATE_4cb8_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2958_l2974_l2963_DUPLICATE_e2fc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2958_l2974_l2963_DUPLICATE_e2fc_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2958_l2974_l2963_l2979_DUPLICATE_b1c1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2958_l2974_l2963_l2979_DUPLICATE_b1c1_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l2969_c30_056c] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_ins;
     sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_x;
     sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_return_output := sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2958_c6_0764] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_left;
     BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output := BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2974_l2963_l2979_l2966_DUPLICATE_ba35 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2974_l2963_l2979_l2966_DUPLICATE_ba35_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2974_c11_5c5e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2974_c7_a7ab] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2974_c7_a7ab_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2979_c11_a26a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2963_c11_afb7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_left;
     BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_return_output := BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2958_l2974_l2963_DUPLICATE_7517 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2958_l2974_l2963_DUPLICATE_7517_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2958_c2_de38_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c6_0764_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2963_c7_6c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2963_c11_afb7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2966_c11_1428_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_5c5e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2979_c11_a26a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2958_l2963_l2966_DUPLICATE_4cb8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2958_l2963_l2966_DUPLICATE_4cb8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2958_l2963_l2966_DUPLICATE_4cb8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2974_l2963_l2979_l2966_DUPLICATE_ba35_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2974_l2963_l2979_l2966_DUPLICATE_ba35_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2974_l2963_l2979_l2966_DUPLICATE_ba35_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2974_l2963_l2979_l2966_DUPLICATE_ba35_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2958_l2974_l2963_DUPLICATE_7517_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2958_l2974_l2963_DUPLICATE_7517_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2958_l2974_l2963_DUPLICATE_7517_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2958_l2974_l2963_l2979_DUPLICATE_b1c1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2958_l2974_l2963_l2979_DUPLICATE_b1c1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2958_l2974_l2963_l2979_DUPLICATE_b1c1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2958_l2974_l2963_l2979_DUPLICATE_b1c1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2958_l2974_l2963_DUPLICATE_e2fc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2958_l2974_l2963_DUPLICATE_e2fc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2958_l2974_l2963_DUPLICATE_e2fc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2974_c7_a7ab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2969_c30_056c_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2974_c7_a7ab] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output := result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2966_c7_c3b2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2974_c7_a7ab] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2979_c7_fd5f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output;

     -- t8_MUX[uxn_opcodes_h_l2966_c7_c3b2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond <= VAR_t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond;
     t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue;
     t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output := t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2958_c1_f670] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2974_c7_a7ab] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2979_c7_fd5f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2959_c3_147d_uxn_opcodes_h_l2959_c3_147d_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2958_c1_f670_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2979_c7_fd5f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2966_c7_c3b2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2966_c7_c3b2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2966_c7_c3b2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2963_c7_6c80] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2974_c7_a7ab] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output;

     -- printf_uxn_opcodes_h_l2959_c3_147d[uxn_opcodes_h_l2959_c3_147d] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2959_c3_147d_uxn_opcodes_h_l2959_c3_147d_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2959_c3_147d_uxn_opcodes_h_l2959_c3_147d_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- t8_MUX[uxn_opcodes_h_l2963_c7_6c80] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2963_c7_6c80_cond <= VAR_t8_MUX_uxn_opcodes_h_l2963_c7_6c80_cond;
     t8_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue;
     t8_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output := t8_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2974_c7_a7ab] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_a7ab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2963_c7_6c80] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output := result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2966_c7_c3b2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2958_c2_de38] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output;

     -- t8_MUX[uxn_opcodes_h_l2958_c2_de38] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2958_c2_de38_cond <= VAR_t8_MUX_uxn_opcodes_h_l2958_c2_de38_cond;
     t8_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue;
     t8_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2958_c2_de38_return_output := t8_MUX_uxn_opcodes_h_l2958_c2_de38_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2963_c7_6c80] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2966_c7_c3b2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2963_c7_6c80] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2966_c7_c3b2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2958_c2_de38_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2958_c2_de38] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_return_output := result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2958_c2_de38] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2958_c2_de38] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2963_c7_6c80] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2963_c7_6c80] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2963_c7_6c80_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2958_c2_de38] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2958_c2_de38] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2984_l2954_DUPLICATE_e679 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2984_l2954_DUPLICATE_e679_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_641b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c2_de38_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c2_de38_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c2_de38_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c2_de38_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c2_de38_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2984_l2954_DUPLICATE_e679_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2984_l2954_DUPLICATE_e679_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
