-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity eor_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor_0CLK_bacf6a1d;
architecture arch of eor_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1035_c6_1e90]
signal BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1035_c1_d6ee]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1035_c2_8def]
signal n8_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1035_c2_8def]
signal t8_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1035_c2_8def]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1035_c2_8def]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1035_c2_8def]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1035_c2_8def]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1035_c2_8def]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1035_c2_8def]
signal result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1036_c3_d954[uxn_opcodes_h_l1036_c3_d954]
signal printf_uxn_opcodes_h_l1036_c3_d954_uxn_opcodes_h_l1036_c3_d954_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1040_c11_75a8]
signal BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1040_c7_bf65]
signal n8_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1040_c7_bf65]
signal t8_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1040_c7_bf65]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1040_c7_bf65]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1040_c7_bf65]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1040_c7_bf65]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1040_c7_bf65]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1040_c7_bf65]
signal result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1043_c11_0d59]
signal BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1043_c7_01fa]
signal n8_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1043_c7_01fa]
signal t8_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1043_c7_01fa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1043_c7_01fa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1043_c7_01fa]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1043_c7_01fa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1043_c7_01fa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1043_c7_01fa]
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1046_c11_d344]
signal BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1046_c7_bb52]
signal n8_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1046_c7_bb52]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1046_c7_bb52]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1046_c7_bb52]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1046_c7_bb52]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1046_c7_bb52]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1046_c7_bb52]
signal result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1049_c30_70cd]
signal sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_return_output : signed(3 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1052_c21_947a]
signal BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_left : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_right : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1054_c11_92d4]
signal BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1054_c7_719b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1054_c7_719b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1054_c7_719b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5b93( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90
BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_left,
BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_right,
BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_return_output);

-- n8_MUX_uxn_opcodes_h_l1035_c2_8def
n8_MUX_uxn_opcodes_h_l1035_c2_8def : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1035_c2_8def_cond,
n8_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue,
n8_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse,
n8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output);

-- t8_MUX_uxn_opcodes_h_l1035_c2_8def
t8_MUX_uxn_opcodes_h_l1035_c2_8def : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1035_c2_8def_cond,
t8_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue,
t8_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse,
t8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_cond,
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_return_output);

-- printf_uxn_opcodes_h_l1036_c3_d954_uxn_opcodes_h_l1036_c3_d954
printf_uxn_opcodes_h_l1036_c3_d954_uxn_opcodes_h_l1036_c3_d954 : entity work.printf_uxn_opcodes_h_l1036_c3_d954_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1036_c3_d954_uxn_opcodes_h_l1036_c3_d954_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8
BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_left,
BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_right,
BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output);

-- n8_MUX_uxn_opcodes_h_l1040_c7_bf65
n8_MUX_uxn_opcodes_h_l1040_c7_bf65 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1040_c7_bf65_cond,
n8_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue,
n8_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse,
n8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output);

-- t8_MUX_uxn_opcodes_h_l1040_c7_bf65
t8_MUX_uxn_opcodes_h_l1040_c7_bf65 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1040_c7_bf65_cond,
t8_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue,
t8_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse,
t8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_cond,
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59
BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_left,
BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_right,
BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output);

-- n8_MUX_uxn_opcodes_h_l1043_c7_01fa
n8_MUX_uxn_opcodes_h_l1043_c7_01fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1043_c7_01fa_cond,
n8_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue,
n8_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse,
n8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output);

-- t8_MUX_uxn_opcodes_h_l1043_c7_01fa
t8_MUX_uxn_opcodes_h_l1043_c7_01fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1043_c7_01fa_cond,
t8_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue,
t8_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse,
t8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_cond,
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344
BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_left,
BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_right,
BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_return_output);

-- n8_MUX_uxn_opcodes_h_l1046_c7_bb52
n8_MUX_uxn_opcodes_h_l1046_c7_bb52 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1046_c7_bb52_cond,
n8_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue,
n8_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse,
n8_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_cond,
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd
sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_ins,
sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_x,
sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_y,
sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a
BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_left,
BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_right,
BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4
BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_left,
BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_right,
BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_return_output,
 n8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output,
 t8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output,
 n8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output,
 t8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output,
 n8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output,
 t8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_return_output,
 n8_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output,
 sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1037_c3_e28e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1036_c3_d954_uxn_opcodes_h_l1036_c3_d954_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1041_c3_642f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1051_c3_a672 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3834_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_9b2d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_d9f7_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_f581_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_29a6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_eeb4_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1060_l1031_DUPLICATE_c7e5_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1051_c3_a672 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1051_c3_a672;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1037_c3_e28e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1037_c3_e28e;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_y := resize(to_signed(-1, 2), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1041_c3_642f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1041_c3_642f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_right := to_unsigned(3, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1054_c11_92d4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1043_c11_0d59] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_left;
     BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output := BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_eeb4 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_eeb4_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1040_c11_75a8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1046_c11_d344] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_left;
     BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_return_output := BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1035_c6_1e90] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_left;
     BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output := BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output;

     -- BIN_OP_XOR[uxn_opcodes_h_l1052_c21_947a] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_left;
     BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_return_output := BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_f581 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_f581_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l1049_c30_70cd] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_ins;
     sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_x;
     sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_return_output := sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_9b2d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_9b2d_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_29a6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_29a6_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3834 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3834_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_d9f7 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_d9f7_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1035_c2_8def_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1035_c2_8def_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_1e90_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1040_c7_bf65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1040_c7_bf65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_75a8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1043_c7_01fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1043_c7_01fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_0d59_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1046_c7_bb52_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_d344_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_92d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_947a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_d9f7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_d9f7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_d9f7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_d9f7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_29a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_29a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_29a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_29a6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_9b2d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_9b2d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_9b2d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_9b2d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3834_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3834_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3834_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3834_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_eeb4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_eeb4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_f581_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_f581_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_f581_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_f581_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_70cd_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1054_c7_719b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_return_output;

     -- n8_MUX[uxn_opcodes_h_l1046_c7_bb52] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1046_c7_bb52_cond <= VAR_n8_MUX_uxn_opcodes_h_l1046_c7_bb52_cond;
     n8_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue;
     n8_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output := n8_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1046_c7_bb52] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;

     -- t8_MUX[uxn_opcodes_h_l1043_c7_01fa] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1043_c7_01fa_cond <= VAR_t8_MUX_uxn_opcodes_h_l1043_c7_01fa_cond;
     t8_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue;
     t8_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output := t8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1046_c7_bb52] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output := result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1046_c7_bb52] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1054_c7_719b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1054_c7_719b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1035_c1_d6ee] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l1036_c3_d954_uxn_opcodes_h_l1036_c3_d954_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_d6ee_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_719b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_719b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_719b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1043_c7_01fa] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output := result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1043_c7_01fa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;

     -- t8_MUX[uxn_opcodes_h_l1040_c7_bf65] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1040_c7_bf65_cond <= VAR_t8_MUX_uxn_opcodes_h_l1040_c7_bf65_cond;
     t8_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue;
     t8_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output := t8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1046_c7_bb52] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;

     -- printf_uxn_opcodes_h_l1036_c3_d954[uxn_opcodes_h_l1036_c3_d954] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1036_c3_d954_uxn_opcodes_h_l1036_c3_d954_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1036_c3_d954_uxn_opcodes_h_l1036_c3_d954_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- n8_MUX[uxn_opcodes_h_l1043_c7_01fa] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1043_c7_01fa_cond <= VAR_n8_MUX_uxn_opcodes_h_l1043_c7_01fa_cond;
     n8_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue;
     n8_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output := n8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1046_c7_bb52] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1046_c7_bb52] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1043_c7_01fa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_bb52_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1043_c7_01fa] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1043_c7_01fa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1040_c7_bf65] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;

     -- n8_MUX[uxn_opcodes_h_l1040_c7_bf65] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1040_c7_bf65_cond <= VAR_n8_MUX_uxn_opcodes_h_l1040_c7_bf65_cond;
     n8_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue;
     n8_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output := n8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;

     -- t8_MUX[uxn_opcodes_h_l1035_c2_8def] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1035_c2_8def_cond <= VAR_t8_MUX_uxn_opcodes_h_l1035_c2_8def_cond;
     t8_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue;
     t8_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output := t8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1040_c7_bf65] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1043_c7_01fa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1040_c7_bf65] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output := result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_01fa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1040_c7_bf65] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1035_c2_8def] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_return_output := result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1035_c2_8def] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_return_output;

     -- n8_MUX[uxn_opcodes_h_l1035_c2_8def] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1035_c2_8def_cond <= VAR_n8_MUX_uxn_opcodes_h_l1035_c2_8def_cond;
     n8_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue;
     n8_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output := n8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1040_c7_bf65] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1035_c2_8def] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1040_c7_bf65] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1035_c2_8def_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_bf65_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1035_c2_8def] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1035_c2_8def] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1035_c2_8def] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1060_l1031_DUPLICATE_c7e5 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1060_l1031_DUPLICATE_c7e5_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5b93(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_8def_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_8def_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_8def_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_8def_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_8def_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1060_l1031_DUPLICATE_c7e5_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1060_l1031_DUPLICATE_c7e5_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
