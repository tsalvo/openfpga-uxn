-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity sub_0CLK_6be78140 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub_0CLK_6be78140;
architecture arch of sub_0CLK_6be78140 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2425_c6_8f21]
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2425_c2_4b4a]
signal n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2425_c2_4b4a]
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2425_c2_4b4a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2425_c2_4b4a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2425_c2_4b4a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2425_c2_4b4a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2425_c2_4b4a]
signal t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2432_c11_5d5e]
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2432_c7_7f6e]
signal n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2432_c7_7f6e]
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2432_c7_7f6e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2432_c7_7f6e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2432_c7_7f6e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2432_c7_7f6e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2432_c7_7f6e]
signal t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2435_c11_a4f9]
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2435_c7_dcb5]
signal n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2435_c7_dcb5]
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2435_c7_dcb5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2435_c7_dcb5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2435_c7_dcb5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2435_c7_dcb5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2435_c7_dcb5]
signal t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2438_c11_fd97]
signal BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2438_c7_7251]
signal n8_MUX_uxn_opcodes_h_l2438_c7_7251_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2438_c7_7251_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2438_c7_7251]
signal result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2438_c7_7251]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2438_c7_7251]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2438_c7_7251]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2438_c7_7251]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2441_c30_67e4]
signal sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_return_output : signed(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2444_c21_fd92]
signal BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2446_c11_2970]
signal BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2446_c7_7280]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2446_c7_7280]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2446_c7_7280]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_return_output : signed(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21
BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_left,
BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_right,
BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_return_output);

-- n8_MUX_uxn_opcodes_h_l2425_c2_4b4a
n8_MUX_uxn_opcodes_h_l2425_c2_4b4a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond,
n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue,
n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse,
n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a
result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output);

-- t8_MUX_uxn_opcodes_h_l2425_c2_4b4a
t8_MUX_uxn_opcodes_h_l2425_c2_4b4a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond,
t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue,
t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse,
t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_left,
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_right,
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_return_output);

-- n8_MUX_uxn_opcodes_h_l2432_c7_7f6e
n8_MUX_uxn_opcodes_h_l2432_c7_7f6e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond,
n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue,
n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse,
n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output);

-- t8_MUX_uxn_opcodes_h_l2432_c7_7f6e
t8_MUX_uxn_opcodes_h_l2432_c7_7f6e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond,
t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue,
t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse,
t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_left,
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_right,
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_return_output);

-- n8_MUX_uxn_opcodes_h_l2435_c7_dcb5
n8_MUX_uxn_opcodes_h_l2435_c7_dcb5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond,
n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue,
n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse,
n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output);

-- t8_MUX_uxn_opcodes_h_l2435_c7_dcb5
t8_MUX_uxn_opcodes_h_l2435_c7_dcb5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond,
t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue,
t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse,
t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97
BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_left,
BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_right,
BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_return_output);

-- n8_MUX_uxn_opcodes_h_l2438_c7_7251
n8_MUX_uxn_opcodes_h_l2438_c7_7251 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2438_c7_7251_cond,
n8_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue,
n8_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse,
n8_MUX_uxn_opcodes_h_l2438_c7_7251_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251
result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_cond,
result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251
result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251
result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251
result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4
sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_ins,
sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_x,
sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_y,
sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92
BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_left,
BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_right,
BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970
BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_left,
BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_right,
BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280
result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280
result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280
result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_return_output,
 n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output,
 t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_return_output,
 n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output,
 t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_return_output,
 n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output,
 t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_return_output,
 n8_MUX_uxn_opcodes_h_l2438_c7_7251_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_return_output,
 sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_ebbb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_ae17 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2438_c7_7251_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2438_c7_7251_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2443_c3_71a8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2447_c3_ac94 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2425_l2438_l2432_l2435_DUPLICATE_cf29_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_7219_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_f68d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2432_l2446_l2435_DUPLICATE_133f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2438_l2435_DUPLICATE_ebd3_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2452_l2421_DUPLICATE_f19e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_ebbb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_ebbb;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2443_c3_71a8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2443_c3_71a8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_ae17 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_ae17;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_right := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2447_c3_ac94 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2447_c3_ac94;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2435_c11_a4f9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2425_l2438_l2432_l2435_DUPLICATE_cf29 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2425_l2438_l2432_l2435_DUPLICATE_cf29_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2432_l2446_l2435_DUPLICATE_133f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2432_l2446_l2435_DUPLICATE_133f_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_f68d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_f68d_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2432_c11_5d5e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2446_c11_2970] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_left;
     BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_return_output := BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2425_c6_8f21] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_left;
     BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_return_output := BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_7219 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_7219_return_output := result.is_stack_write;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2444_c21_fd92] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2438_c11_fd97] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_left;
     BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_return_output := BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2441_c30_67e4] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_ins;
     sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_x;
     sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_return_output := sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2438_l2435_DUPLICATE_ebd3 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2438_l2435_DUPLICATE_ebd3_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c6_8f21_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_5d5e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_a4f9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2438_c7_7251_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_fd97_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2446_c11_2970_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2444_c21_fd92_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_f68d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_f68d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_f68d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_f68d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2432_l2446_l2435_DUPLICATE_133f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2432_l2446_l2435_DUPLICATE_133f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2432_l2446_l2435_DUPLICATE_133f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2432_l2446_l2435_DUPLICATE_133f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_7219_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_7219_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_7219_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2425_l2432_l2446_l2435_DUPLICATE_7219_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2438_l2435_DUPLICATE_ebd3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2438_l2435_DUPLICATE_ebd3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2425_l2438_l2432_l2435_DUPLICATE_cf29_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2425_l2438_l2432_l2435_DUPLICATE_cf29_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2425_l2438_l2432_l2435_DUPLICATE_cf29_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2425_l2438_l2432_l2435_DUPLICATE_cf29_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2441_c30_67e4_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2446_c7_7280] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2446_c7_7280] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2438_c7_7251] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2446_c7_7280] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_return_output;

     -- t8_MUX[uxn_opcodes_h_l2435_c7_dcb5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond <= VAR_t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond;
     t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue;
     t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output := t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2438_c7_7251] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_return_output := result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_return_output;

     -- n8_MUX[uxn_opcodes_h_l2438_c7_7251] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2438_c7_7251_cond <= VAR_n8_MUX_uxn_opcodes_h_l2438_c7_7251_cond;
     n8_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue;
     n8_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2438_c7_7251_return_output := n8_MUX_uxn_opcodes_h_l2438_c7_7251_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2438_c7_7251_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2446_c7_7280_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2446_c7_7280_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2446_c7_7280_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2438_c7_7251_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2438_c7_7251_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2438_c7_7251] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2435_c7_dcb5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output := result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2435_c7_dcb5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2438_c7_7251] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_return_output;

     -- t8_MUX[uxn_opcodes_h_l2432_c7_7f6e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond <= VAR_t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond;
     t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue;
     t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output := t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2435_c7_dcb5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond <= VAR_n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond;
     n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue;
     n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output := n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2438_c7_7251] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_7251_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_7251_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2438_c7_7251_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2432_c7_7f6e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2435_c7_dcb5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;

     -- t8_MUX[uxn_opcodes_h_l2425_c2_4b4a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond <= VAR_t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond;
     t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue;
     t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output := t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output;

     -- n8_MUX[uxn_opcodes_h_l2432_c7_7f6e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond <= VAR_n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond;
     n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue;
     n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output := n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2432_c7_7f6e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2435_c7_dcb5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2435_c7_dcb5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_dcb5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2432_c7_7f6e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2425_c2_4b4a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2425_c2_4b4a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2432_c7_7f6e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2432_c7_7f6e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2425_c2_4b4a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond <= VAR_n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond;
     n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue;
     n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output := n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_7f6e_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2425_c2_4b4a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2425_c2_4b4a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2425_c2_4b4a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2452_l2421_DUPLICATE_f19e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2452_l2421_DUPLICATE_f19e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c2_4b4a_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2452_l2421_DUPLICATE_f19e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2452_l2421_DUPLICATE_f19e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
