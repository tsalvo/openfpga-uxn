-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity ora_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ora_0CLK_bacf6a1d;
architecture arch of ora_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l956_c6_8616]
signal BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l956_c1_f73c]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l956_c2_b257]
signal t8_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l956_c2_b257]
signal n8_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l956_c2_b257]
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l956_c2_b257]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l956_c2_b257]
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l956_c2_b257]
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l956_c2_b257]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l956_c2_b257]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l957_c3_4c98[uxn_opcodes_h_l957_c3_4c98]
signal printf_uxn_opcodes_h_l957_c3_4c98_uxn_opcodes_h_l957_c3_4c98_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l961_c11_8d42]
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l961_c7_c022]
signal t8_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l961_c7_c022]
signal n8_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l961_c7_c022]
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l961_c7_c022]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l961_c7_c022]
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l961_c7_c022]
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l961_c7_c022]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l961_c7_c022]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l964_c11_65db]
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l964_c7_b68b]
signal t8_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l964_c7_b68b]
signal n8_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l964_c7_b68b]
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l964_c7_b68b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l964_c7_b68b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l964_c7_b68b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l964_c7_b68b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l964_c7_b68b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l967_c11_a6f9]
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l967_c7_bb45]
signal n8_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l967_c7_bb45]
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l967_c7_bb45]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l967_c7_bb45]
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l967_c7_bb45]
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l967_c7_bb45]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l967_c7_bb45]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l970_c30_dbcf]
signal sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l973_c21_64c7]
signal BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_left : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_right : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l975_c11_d5dd]
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l975_c7_9ac6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l975_c7_9ac6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l975_c7_9ac6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616
BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_left,
BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_right,
BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_return_output);

-- t8_MUX_uxn_opcodes_h_l956_c2_b257
t8_MUX_uxn_opcodes_h_l956_c2_b257 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l956_c2_b257_cond,
t8_MUX_uxn_opcodes_h_l956_c2_b257_iftrue,
t8_MUX_uxn_opcodes_h_l956_c2_b257_iffalse,
t8_MUX_uxn_opcodes_h_l956_c2_b257_return_output);

-- n8_MUX_uxn_opcodes_h_l956_c2_b257
n8_MUX_uxn_opcodes_h_l956_c2_b257 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l956_c2_b257_cond,
n8_MUX_uxn_opcodes_h_l956_c2_b257_iftrue,
n8_MUX_uxn_opcodes_h_l956_c2_b257_iffalse,
n8_MUX_uxn_opcodes_h_l956_c2_b257_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257
result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_cond,
result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output);

-- printf_uxn_opcodes_h_l957_c3_4c98_uxn_opcodes_h_l957_c3_4c98
printf_uxn_opcodes_h_l957_c3_4c98_uxn_opcodes_h_l957_c3_4c98 : entity work.printf_uxn_opcodes_h_l957_c3_4c98_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l957_c3_4c98_uxn_opcodes_h_l957_c3_4c98_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42
BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_left,
BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_right,
BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output);

-- t8_MUX_uxn_opcodes_h_l961_c7_c022
t8_MUX_uxn_opcodes_h_l961_c7_c022 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l961_c7_c022_cond,
t8_MUX_uxn_opcodes_h_l961_c7_c022_iftrue,
t8_MUX_uxn_opcodes_h_l961_c7_c022_iffalse,
t8_MUX_uxn_opcodes_h_l961_c7_c022_return_output);

-- n8_MUX_uxn_opcodes_h_l961_c7_c022
n8_MUX_uxn_opcodes_h_l961_c7_c022 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l961_c7_c022_cond,
n8_MUX_uxn_opcodes_h_l961_c7_c022_iftrue,
n8_MUX_uxn_opcodes_h_l961_c7_c022_iffalse,
n8_MUX_uxn_opcodes_h_l961_c7_c022_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022
result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_cond,
result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db
BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_left,
BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_right,
BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output);

-- t8_MUX_uxn_opcodes_h_l964_c7_b68b
t8_MUX_uxn_opcodes_h_l964_c7_b68b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l964_c7_b68b_cond,
t8_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue,
t8_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse,
t8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output);

-- n8_MUX_uxn_opcodes_h_l964_c7_b68b
n8_MUX_uxn_opcodes_h_l964_c7_b68b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l964_c7_b68b_cond,
n8_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue,
n8_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse,
n8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b
result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_cond,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9
BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_left,
BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_right,
BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_return_output);

-- n8_MUX_uxn_opcodes_h_l967_c7_bb45
n8_MUX_uxn_opcodes_h_l967_c7_bb45 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l967_c7_bb45_cond,
n8_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue,
n8_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse,
n8_MUX_uxn_opcodes_h_l967_c7_bb45_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45
result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_cond,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output);

-- sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf
sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_ins,
sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_x,
sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_y,
sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7
BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7 : entity work.BIN_OP_OR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_left,
BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_right,
BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd
BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_left,
BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_right,
BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_return_output,
 t8_MUX_uxn_opcodes_h_l956_c2_b257_return_output,
 n8_MUX_uxn_opcodes_h_l956_c2_b257_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output,
 t8_MUX_uxn_opcodes_h_l961_c7_c022_return_output,
 n8_MUX_uxn_opcodes_h_l961_c7_c022_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output,
 t8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output,
 n8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_return_output,
 n8_MUX_uxn_opcodes_h_l967_c7_bb45_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output,
 sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_return_output,
 BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_fbb6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l957_c3_4c98_uxn_opcodes_h_l957_c3_4c98_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_dc29 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_43cd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_9969_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_c727_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_1190_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_64fc_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l964_l967_l961_l975_DUPLICATE_6dbd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_dd3a_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l981_l952_DUPLICATE_b498_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_fbb6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_fbb6;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_right := to_unsigned(4, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_43cd := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_43cd;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_dc29 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_dc29;
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_b257_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_c022_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_b257_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_c022_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l961_c11_8d42] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_left;
     BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output := BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_c727 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_c727_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_1190 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_1190_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_9969 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_9969_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l956_c6_8616] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_left;
     BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output := BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_dd3a LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_dd3a_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_64fc LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_64fc_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l964_c11_65db] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_left;
     BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output := BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l975_c11_d5dd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_left;
     BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_return_output := BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l973_c21_64c7] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_left;
     BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_return_output := BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l964_l967_l961_l975_DUPLICATE_6dbd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l964_l967_l961_l975_DUPLICATE_6dbd_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l970_c30_dbcf] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_ins;
     sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_x <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_x;
     sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_y <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_return_output := sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l967_c11_a6f9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_left;
     BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_return_output := BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_b257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_b257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_8616_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_c022_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_c022_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_8d42_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_b68b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_b68b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_65db_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_bb45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_a6f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_d5dd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_64c7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_64fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_64fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_64fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_64fc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l964_l967_l961_l975_DUPLICATE_6dbd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l964_l967_l961_l975_DUPLICATE_6dbd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l964_l967_l961_l975_DUPLICATE_6dbd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l964_l967_l961_l975_DUPLICATE_6dbd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_c727_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_c727_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_c727_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_c727_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_1190_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_1190_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_1190_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l964_l956_l961_l975_DUPLICATE_1190_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_dd3a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l964_l967_DUPLICATE_dd3a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_9969_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_9969_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_9969_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l964_l956_l967_l961_DUPLICATE_9969_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_dbcf_return_output;
     -- n8_MUX[uxn_opcodes_h_l967_c7_bb45] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l967_c7_bb45_cond <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_bb45_cond;
     n8_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue;
     n8_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_bb45_return_output := n8_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l967_c7_bb45] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l975_c7_9ac6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l956_c1_f73c] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l975_c7_9ac6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output;

     -- t8_MUX[uxn_opcodes_h_l964_c7_b68b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l964_c7_b68b_cond <= VAR_t8_MUX_uxn_opcodes_h_l964_c7_b68b_cond;
     t8_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue;
     t8_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output := t8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l967_c7_bb45] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_cond;
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_return_output := result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l975_c7_9ac6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l967_c7_bb45] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l957_c3_4c98_uxn_opcodes_h_l957_c3_4c98_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_f73c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_9ac6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_c022_iffalse := VAR_t8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l967_c7_bb45] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l964_c7_b68b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_return_output := result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;

     -- n8_MUX[uxn_opcodes_h_l964_c7_b68b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l964_c7_b68b_cond <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_b68b_cond;
     n8_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue;
     n8_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output := n8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l964_c7_b68b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;

     -- printf_uxn_opcodes_h_l957_c3_4c98[uxn_opcodes_h_l957_c3_4c98] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l957_c3_4c98_uxn_opcodes_h_l957_c3_4c98_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l957_c3_4c98_uxn_opcodes_h_l957_c3_4c98_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l964_c7_b68b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l967_c7_bb45] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l967_c7_bb45] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;

     -- t8_MUX[uxn_opcodes_h_l961_c7_c022] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l961_c7_c022_cond <= VAR_t8_MUX_uxn_opcodes_h_l961_c7_c022_cond;
     t8_MUX_uxn_opcodes_h_l961_c7_c022_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l961_c7_c022_iftrue;
     t8_MUX_uxn_opcodes_h_l961_c7_c022_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l961_c7_c022_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_c022_return_output := t8_MUX_uxn_opcodes_h_l961_c7_c022_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_c022_iffalse := VAR_n8_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_bb45_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_b257_iffalse := VAR_t8_MUX_uxn_opcodes_h_l961_c7_c022_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l964_c7_b68b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l961_c7_c022] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_cond;
     result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_return_output := result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l961_c7_c022] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l964_c7_b68b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;

     -- n8_MUX[uxn_opcodes_h_l961_c7_c022] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l961_c7_c022_cond <= VAR_n8_MUX_uxn_opcodes_h_l961_c7_c022_cond;
     n8_MUX_uxn_opcodes_h_l961_c7_c022_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l961_c7_c022_iftrue;
     n8_MUX_uxn_opcodes_h_l961_c7_c022_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l961_c7_c022_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_c022_return_output := n8_MUX_uxn_opcodes_h_l961_c7_c022_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l964_c7_b68b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;

     -- t8_MUX[uxn_opcodes_h_l956_c2_b257] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l956_c2_b257_cond <= VAR_t8_MUX_uxn_opcodes_h_l956_c2_b257_cond;
     t8_MUX_uxn_opcodes_h_l956_c2_b257_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l956_c2_b257_iftrue;
     t8_MUX_uxn_opcodes_h_l956_c2_b257_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l956_c2_b257_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_b257_return_output := t8_MUX_uxn_opcodes_h_l956_c2_b257_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l961_c7_c022] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_b257_iffalse := VAR_n8_MUX_uxn_opcodes_h_l961_c7_c022_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_b68b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_c022_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_c022_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l956_c2_b257_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l961_c7_c022] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l961_c7_c022] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l956_c2_b257] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_cond;
     result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_return_output := result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l961_c7_c022] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l956_c2_b257] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l956_c2_b257] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output;

     -- n8_MUX[uxn_opcodes_h_l956_c2_b257] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l956_c2_b257_cond <= VAR_n8_MUX_uxn_opcodes_h_l956_c2_b257_cond;
     n8_MUX_uxn_opcodes_h_l956_c2_b257_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l956_c2_b257_iftrue;
     n8_MUX_uxn_opcodes_h_l956_c2_b257_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l956_c2_b257_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_b257_return_output := n8_MUX_uxn_opcodes_h_l956_c2_b257_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l956_c2_b257_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_c022_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_c022_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_c022_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l956_c2_b257] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l956_c2_b257] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l956_c2_b257] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l981_l952_DUPLICATE_b498 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l981_l952_DUPLICATE_b498_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_b257_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_b257_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_b257_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_b257_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_b257_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l981_l952_DUPLICATE_b498_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l981_l952_DUPLICATE_b498_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
