-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity str1_0CLK_faaf4b1a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end str1_0CLK_faaf4b1a;
architecture arch of str1_0CLK_faaf4b1a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1596_c6_4ff0]
signal BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1596_c1_4631]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1596_c2_1595]
signal n8_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1596_c2_1595]
signal t8_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1596_c2_1595]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1596_c2_1595]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1596_c2_1595]
signal result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1596_c2_1595]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1596_c2_1595]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1596_c2_1595]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1596_c2_1595]
signal result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l1597_c3_b2bf[uxn_opcodes_h_l1597_c3_b2bf]
signal printf_uxn_opcodes_h_l1597_c3_b2bf_uxn_opcodes_h_l1597_c3_b2bf_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1601_c11_e799]
signal BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1601_c7_d453]
signal n8_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1601_c7_d453]
signal t8_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1601_c7_d453]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1601_c7_d453]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1601_c7_d453]
signal result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1601_c7_d453]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1601_c7_d453]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1601_c7_d453]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1601_c7_d453]
signal result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1604_c11_ce14]
signal BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1604_c7_f6d0]
signal n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1604_c7_f6d0]
signal t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1604_c7_f6d0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1604_c7_f6d0]
signal result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1604_c7_f6d0]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1604_c7_f6d0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1604_c7_f6d0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1604_c7_f6d0]
signal result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1607_c11_757e]
signal BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1607_c7_38a0]
signal n8_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1607_c7_38a0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1607_c7_38a0]
signal result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1607_c7_38a0]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1607_c7_38a0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1607_c7_38a0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1607_c7_38a0]
signal result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1610_c30_11d7]
signal sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1612_c22_dde5]
signal BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1615_c11_ea83]
signal BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1615_c7_9e06]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1615_c7_9e06]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1615_c7_9e06]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_18d1( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : signed;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.sp_relative_shift := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_sp_shift := ref_toks_6;
      base.u16_value := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0
BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_left,
BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_right,
BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_return_output);

-- n8_MUX_uxn_opcodes_h_l1596_c2_1595
n8_MUX_uxn_opcodes_h_l1596_c2_1595 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1596_c2_1595_cond,
n8_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue,
n8_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse,
n8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output);

-- t8_MUX_uxn_opcodes_h_l1596_c2_1595
t8_MUX_uxn_opcodes_h_l1596_c2_1595 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1596_c2_1595_cond,
t8_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue,
t8_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse,
t8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595
result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595
result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_cond,
result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595
result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595
result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595
result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595
result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_cond,
result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output);

-- printf_uxn_opcodes_h_l1597_c3_b2bf_uxn_opcodes_h_l1597_c3_b2bf
printf_uxn_opcodes_h_l1597_c3_b2bf_uxn_opcodes_h_l1597_c3_b2bf : entity work.printf_uxn_opcodes_h_l1597_c3_b2bf_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1597_c3_b2bf_uxn_opcodes_h_l1597_c3_b2bf_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799
BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_left,
BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_right,
BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output);

-- n8_MUX_uxn_opcodes_h_l1601_c7_d453
n8_MUX_uxn_opcodes_h_l1601_c7_d453 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1601_c7_d453_cond,
n8_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue,
n8_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse,
n8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output);

-- t8_MUX_uxn_opcodes_h_l1601_c7_d453
t8_MUX_uxn_opcodes_h_l1601_c7_d453 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1601_c7_d453_cond,
t8_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue,
t8_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse,
t8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453
result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453
result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_cond,
result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453
result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453
result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453
result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453
result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_cond,
result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14
BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_left,
BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_right,
BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output);

-- n8_MUX_uxn_opcodes_h_l1604_c7_f6d0
n8_MUX_uxn_opcodes_h_l1604_c7_f6d0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond,
n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue,
n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse,
n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output);

-- t8_MUX_uxn_opcodes_h_l1604_c7_f6d0
t8_MUX_uxn_opcodes_h_l1604_c7_f6d0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond,
t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue,
t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse,
t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0
result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0
result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0
result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond,
result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e
BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_left,
BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_right,
BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_return_output);

-- n8_MUX_uxn_opcodes_h_l1607_c7_38a0
n8_MUX_uxn_opcodes_h_l1607_c7_38a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1607_c7_38a0_cond,
n8_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue,
n8_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse,
n8_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0
result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0
result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0
result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0
result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0
result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_cond,
result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7
sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_ins,
sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_x,
sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_y,
sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5
BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_left,
BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_right,
BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83
BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_left,
BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_right,
BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06
result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06
result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_return_output,
 n8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
 t8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output,
 n8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output,
 t8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output,
 n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output,
 t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_return_output,
 n8_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output,
 sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1598_c3_0002 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1597_c3_b2bf_uxn_opcodes_h_l1597_c3_b2bf_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1602_c3_b9a9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1601_c7_d453_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1612_c3_ae2b : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1612_c27_42f6_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_ba71_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_a722_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_a8d1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_e23b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_682d_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1604_l1607_l1601_DUPLICATE_c6b8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_18d1_uxn_opcodes_h_l1621_l1592_DUPLICATE_0259_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_iffalse := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_right := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_y := resize(to_signed(-2, 3), 4);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1602_c3_b9a9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1602_c3_b9a9;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1598_c3_0002 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1598_c3_0002;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse := n8;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse := t8;
     -- CAST_TO_int8_t[uxn_opcodes_h_l1612_c27_42f6] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1612_c27_42f6_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- sp_relative_shift[uxn_opcodes_h_l1610_c30_11d7] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_ins;
     sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_x;
     sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_return_output := sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_682d LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_682d_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_a8d1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_a8d1_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1596_c6_4ff0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_e23b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_e23b_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1607_c11_757e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1615_c11_ea83] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_left;
     BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_return_output := BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1604_c11_ce14] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_left;
     BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output := BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_ba71 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_ba71_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1601_c11_e799] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_left;
     BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output := BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_a722 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_a722_return_output := result.u8_value;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1601_c7_d453] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1601_c7_d453_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1604_l1607_l1601_DUPLICATE_c6b8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1604_l1607_l1601_DUPLICATE_c6b8_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1596_c2_1595_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1596_c2_1595_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1596_c6_4ff0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1601_c7_d453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1601_c7_d453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_e799_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c11_ce14_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1607_c7_38a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1607_c11_757e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_ea83_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1612_c27_42f6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_ba71_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_ba71_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_ba71_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_ba71_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_682d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_682d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_682d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_682d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1604_l1607_l1601_DUPLICATE_c6b8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1604_l1607_l1601_DUPLICATE_c6b8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1604_l1607_l1601_DUPLICATE_c6b8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1604_l1607_l1601_DUPLICATE_c6b8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_a8d1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_a8d1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_a8d1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_a8d1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_e23b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_e23b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_e23b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1615_l1604_l1596_l1601_DUPLICATE_e23b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_a722_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_a722_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_a722_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1604_l1596_l1607_l1601_DUPLICATE_a722_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1601_c7_d453_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1610_c30_11d7_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1615_c7_9e06] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1615_c7_9e06] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1615_c7_9e06] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output;

     -- t8_MUX[uxn_opcodes_h_l1604_c7_f6d0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond <= VAR_t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond;
     t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue;
     t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output := t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1607_c7_38a0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1607_c7_38a0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1601_c7_d453] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;

     -- n8_MUX[uxn_opcodes_h_l1607_c7_38a0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1607_c7_38a0_cond <= VAR_n8_MUX_uxn_opcodes_h_l1607_c7_38a0_cond;
     n8_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue;
     n8_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output := n8_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1596_c1_4631] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1612_c22_dde5] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1612_c3_ae2b := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1612_c22_dde5_return_output)),16);
     VAR_printf_uxn_opcodes_h_l1597_c3_b2bf_uxn_opcodes_h_l1597_c3_b2bf_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1596_c1_4631_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_9e06_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1612_c3_ae2b;
     -- t8_MUX[uxn_opcodes_h_l1601_c7_d453] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1601_c7_d453_cond <= VAR_t8_MUX_uxn_opcodes_h_l1601_c7_d453_cond;
     t8_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue;
     t8_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output := t8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1596_c2_1595] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1607_c7_38a0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1604_c7_f6d0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1604_c7_f6d0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1607_c7_38a0] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1607_c7_38a0] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output := result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;

     -- printf_uxn_opcodes_h_l1597_c3_b2bf[uxn_opcodes_h_l1597_c3_b2bf] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1597_c3_b2bf_uxn_opcodes_h_l1597_c3_b2bf_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1597_c3_b2bf_uxn_opcodes_h_l1597_c3_b2bf_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- n8_MUX[uxn_opcodes_h_l1604_c7_f6d0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond <= VAR_n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond;
     n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue;
     n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output := n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1607_c7_38a0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1607_c7_38a0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;
     -- n8_MUX[uxn_opcodes_h_l1601_c7_d453] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1601_c7_d453_cond <= VAR_n8_MUX_uxn_opcodes_h_l1601_c7_d453_cond;
     n8_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue;
     n8_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output := n8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1601_c7_d453] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1601_c7_d453] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output := result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1604_c7_f6d0] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1604_c7_f6d0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1604_c7_f6d0] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output := result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;

     -- t8_MUX[uxn_opcodes_h_l1596_c2_1595] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1596_c2_1595_cond <= VAR_t8_MUX_uxn_opcodes_h_l1596_c2_1595_cond;
     t8_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue;
     t8_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output := t8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1604_c7_f6d0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c7_f6d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1596_c2_1595] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1601_c7_d453] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1601_c7_d453] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output := result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1601_c7_d453] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;

     -- n8_MUX[uxn_opcodes_h_l1596_c2_1595] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1596_c2_1595_cond <= VAR_n8_MUX_uxn_opcodes_h_l1596_c2_1595_cond;
     n8_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue;
     n8_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output := n8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1596_c2_1595] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output := result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1601_c7_d453] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1596_c2_1595_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_d453_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1596_c2_1595] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1596_c2_1595] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1596_c2_1595] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output := result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1596_c2_1595] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_18d1_uxn_opcodes_h_l1621_l1592_DUPLICATE_0259 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_18d1_uxn_opcodes_h_l1621_l1592_DUPLICATE_0259_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_18d1(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1596_c2_1595_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1596_c2_1595_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_18d1_uxn_opcodes_h_l1621_l1592_DUPLICATE_0259_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_18d1_uxn_opcodes_h_l1621_l1592_DUPLICATE_0259_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
