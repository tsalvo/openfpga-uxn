-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity add_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end add_0CLK_bacf6a1d;
architecture arch of add_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l798_c6_693d]
signal BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l798_c1_c4e2]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l798_c2_0643]
signal t8_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l798_c2_0643]
signal n8_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l798_c2_0643]
signal result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l798_c2_0643]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l798_c2_0643]
signal result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l798_c2_0643]
signal result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l798_c2_0643]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l798_c2_0643]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l799_c3_e737[uxn_opcodes_h_l799_c3_e737]
signal printf_uxn_opcodes_h_l799_c3_e737_uxn_opcodes_h_l799_c3_e737_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l803_c11_0251]
signal BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l803_c7_90ad]
signal t8_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l803_c7_90ad]
signal n8_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l803_c7_90ad]
signal result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l803_c7_90ad]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l803_c7_90ad]
signal result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l803_c7_90ad]
signal result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l803_c7_90ad]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l803_c7_90ad]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l806_c11_9f10]
signal BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l806_c7_1307]
signal t8_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l806_c7_1307]
signal n8_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l806_c7_1307]
signal result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l806_c7_1307]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l806_c7_1307]
signal result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l806_c7_1307]
signal result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l806_c7_1307]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l806_c7_1307]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l809_c11_7f2b]
signal BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l809_c7_0507]
signal n8_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l809_c7_0507_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l809_c7_0507]
signal result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l809_c7_0507]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l809_c7_0507]
signal result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l809_c7_0507]
signal result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l809_c7_0507]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l809_c7_0507]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l812_c30_942f]
signal sp_relative_shift_uxn_opcodes_h_l812_c30_942f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l812_c30_942f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l812_c30_942f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l812_c30_942f_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l815_c21_79e0]
signal BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_right : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l817_c11_06b4]
signal BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l817_c7_6b33]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l817_c7_6b33]
signal result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l817_c7_6b33]
signal result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d
BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_left,
BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_right,
BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_return_output);

-- t8_MUX_uxn_opcodes_h_l798_c2_0643
t8_MUX_uxn_opcodes_h_l798_c2_0643 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l798_c2_0643_cond,
t8_MUX_uxn_opcodes_h_l798_c2_0643_iftrue,
t8_MUX_uxn_opcodes_h_l798_c2_0643_iffalse,
t8_MUX_uxn_opcodes_h_l798_c2_0643_return_output);

-- n8_MUX_uxn_opcodes_h_l798_c2_0643
n8_MUX_uxn_opcodes_h_l798_c2_0643 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l798_c2_0643_cond,
n8_MUX_uxn_opcodes_h_l798_c2_0643_iftrue,
n8_MUX_uxn_opcodes_h_l798_c2_0643_iffalse,
n8_MUX_uxn_opcodes_h_l798_c2_0643_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643
result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_cond,
result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643
result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643
result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643
result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643
result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output);

-- printf_uxn_opcodes_h_l799_c3_e737_uxn_opcodes_h_l799_c3_e737
printf_uxn_opcodes_h_l799_c3_e737_uxn_opcodes_h_l799_c3_e737 : entity work.printf_uxn_opcodes_h_l799_c3_e737_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l799_c3_e737_uxn_opcodes_h_l799_c3_e737_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251
BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_left,
BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_right,
BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output);

-- t8_MUX_uxn_opcodes_h_l803_c7_90ad
t8_MUX_uxn_opcodes_h_l803_c7_90ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l803_c7_90ad_cond,
t8_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue,
t8_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse,
t8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output);

-- n8_MUX_uxn_opcodes_h_l803_c7_90ad
n8_MUX_uxn_opcodes_h_l803_c7_90ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l803_c7_90ad_cond,
n8_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue,
n8_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse,
n8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad
result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_cond,
result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad
result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad
result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad
result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad
result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10
BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_left,
BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_right,
BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output);

-- t8_MUX_uxn_opcodes_h_l806_c7_1307
t8_MUX_uxn_opcodes_h_l806_c7_1307 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l806_c7_1307_cond,
t8_MUX_uxn_opcodes_h_l806_c7_1307_iftrue,
t8_MUX_uxn_opcodes_h_l806_c7_1307_iffalse,
t8_MUX_uxn_opcodes_h_l806_c7_1307_return_output);

-- n8_MUX_uxn_opcodes_h_l806_c7_1307
n8_MUX_uxn_opcodes_h_l806_c7_1307 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l806_c7_1307_cond,
n8_MUX_uxn_opcodes_h_l806_c7_1307_iftrue,
n8_MUX_uxn_opcodes_h_l806_c7_1307_iffalse,
n8_MUX_uxn_opcodes_h_l806_c7_1307_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307
result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_cond,
result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307
result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307
result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307
result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307
result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b
BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_left,
BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_right,
BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_return_output);

-- n8_MUX_uxn_opcodes_h_l809_c7_0507
n8_MUX_uxn_opcodes_h_l809_c7_0507 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l809_c7_0507_cond,
n8_MUX_uxn_opcodes_h_l809_c7_0507_iftrue,
n8_MUX_uxn_opcodes_h_l809_c7_0507_iffalse,
n8_MUX_uxn_opcodes_h_l809_c7_0507_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507
result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_cond,
result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507
result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507
result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507
result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507
result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output);

-- sp_relative_shift_uxn_opcodes_h_l812_c30_942f
sp_relative_shift_uxn_opcodes_h_l812_c30_942f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l812_c30_942f_ins,
sp_relative_shift_uxn_opcodes_h_l812_c30_942f_x,
sp_relative_shift_uxn_opcodes_h_l812_c30_942f_y,
sp_relative_shift_uxn_opcodes_h_l812_c30_942f_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0
BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0 : entity work.BIN_OP_PLUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_left,
BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_right,
BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4
BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_left,
BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_right,
BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33
result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33
result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33
result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_return_output,
 t8_MUX_uxn_opcodes_h_l798_c2_0643_return_output,
 n8_MUX_uxn_opcodes_h_l798_c2_0643_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output,
 t8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output,
 n8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output,
 t8_MUX_uxn_opcodes_h_l806_c7_1307_return_output,
 n8_MUX_uxn_opcodes_h_l806_c7_1307_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_return_output,
 n8_MUX_uxn_opcodes_h_l809_c7_0507_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output,
 sp_relative_shift_uxn_opcodes_h_l812_c30_942f_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l800_c3_8bbc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l799_c3_e737_uxn_opcodes_h_l799_c3_e737_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l804_c3_acd3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l809_c7_0507_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l815_c3_eda0 : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l814_c3_af57 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l812_c30_942f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l812_c30_942f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l812_c30_942f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l812_c30_942f_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_return_output : unsigned(8 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_def5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_55f8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_098c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_6c55_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l803_l817_l806_l809_DUPLICATE_e8f8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l806_l809_DUPLICATE_b501_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l823_l794_DUPLICATE_89d4_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l812_c30_942f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l804_c3_acd3 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l804_c3_acd3;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l812_c30_942f_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l814_c3_af57 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l814_c3_af57;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l800_c3_8bbc := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l800_c3_8bbc;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l812_c30_942f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l798_c2_0643_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l806_c7_1307_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l809_c7_0507_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l809_c7_0507_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l806_c7_1307_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l798_c2_0643_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l806_c7_1307_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l803_c11_0251] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_left;
     BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output := BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l812_c30_942f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l812_c30_942f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l812_c30_942f_ins;
     sp_relative_shift_uxn_opcodes_h_l812_c30_942f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l812_c30_942f_x;
     sp_relative_shift_uxn_opcodes_h_l812_c30_942f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l812_c30_942f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l812_c30_942f_return_output := sp_relative_shift_uxn_opcodes_h_l812_c30_942f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l806_c11_9f10] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_left;
     BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output := BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_def5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_def5_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_6c55 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_6c55_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l798_c6_693d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_left;
     BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output := BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_098c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_098c_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l803_l817_l806_l809_DUPLICATE_e8f8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l803_l817_l806_l809_DUPLICATE_e8f8_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l806_l809_DUPLICATE_b501 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l806_l809_DUPLICATE_b501_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l809_c11_7f2b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_left;
     BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_return_output := BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l817_c11_06b4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_left;
     BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_return_output := BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l815_c21_79e0] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_left;
     BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_return_output := BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_55f8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_55f8_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l798_c2_0643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l798_c2_0643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l798_c6_693d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l803_c7_90ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l803_c7_90ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l803_c11_0251_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l806_c7_1307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l806_c7_1307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l806_c11_9f10_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l809_c7_0507_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l809_c11_7f2b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l817_c11_06b4_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l815_c3_eda0 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l815_c21_79e0_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_6c55_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_6c55_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_6c55_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_6c55_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l803_l817_l806_l809_DUPLICATE_e8f8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l803_l817_l806_l809_DUPLICATE_e8f8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l803_l817_l806_l809_DUPLICATE_e8f8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l803_l817_l806_l809_DUPLICATE_e8f8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_55f8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_55f8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_55f8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_55f8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_098c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_098c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_098c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l803_l817_l806_l798_DUPLICATE_098c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l806_l809_DUPLICATE_b501_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l806_l809_DUPLICATE_b501_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_def5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_def5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_def5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l803_l806_l798_l809_DUPLICATE_def5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l812_c30_942f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_iftrue := VAR_result_u8_value_uxn_opcodes_h_l815_c3_eda0;
     -- result_u8_value_MUX[uxn_opcodes_h_l809_c7_0507] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_cond;
     result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_return_output := result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_return_output;

     -- n8_MUX[uxn_opcodes_h_l809_c7_0507] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l809_c7_0507_cond <= VAR_n8_MUX_uxn_opcodes_h_l809_c7_0507_cond;
     n8_MUX_uxn_opcodes_h_l809_c7_0507_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l809_c7_0507_iftrue;
     n8_MUX_uxn_opcodes_h_l809_c7_0507_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l809_c7_0507_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l809_c7_0507_return_output := n8_MUX_uxn_opcodes_h_l809_c7_0507_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l798_c1_c4e2] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l817_c7_6b33] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l817_c7_6b33] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l809_c7_0507] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l809_c7_0507] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_return_output;

     -- t8_MUX[uxn_opcodes_h_l806_c7_1307] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l806_c7_1307_cond <= VAR_t8_MUX_uxn_opcodes_h_l806_c7_1307_cond;
     t8_MUX_uxn_opcodes_h_l806_c7_1307_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l806_c7_1307_iftrue;
     t8_MUX_uxn_opcodes_h_l806_c7_1307_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l806_c7_1307_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l806_c7_1307_return_output := t8_MUX_uxn_opcodes_h_l806_c7_1307_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l817_c7_6b33] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l799_c3_e737_uxn_opcodes_h_l799_c3_e737_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l798_c1_c4e2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l806_c7_1307_iffalse := VAR_n8_MUX_uxn_opcodes_h_l809_c7_0507_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l817_c7_6b33_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l817_c7_6b33_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l817_c7_6b33_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l809_c7_0507_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l809_c7_0507_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse := VAR_t8_MUX_uxn_opcodes_h_l806_c7_1307_return_output;
     -- printf_uxn_opcodes_h_l799_c3_e737[uxn_opcodes_h_l799_c3_e737] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l799_c3_e737_uxn_opcodes_h_l799_c3_e737_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l799_c3_e737_uxn_opcodes_h_l799_c3_e737_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_opc_done_MUX[uxn_opcodes_h_l809_c7_0507] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l809_c7_0507] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l806_c7_1307] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l806_c7_1307] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_cond;
     result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_return_output := result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_return_output;

     -- t8_MUX[uxn_opcodes_h_l803_c7_90ad] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l803_c7_90ad_cond <= VAR_t8_MUX_uxn_opcodes_h_l803_c7_90ad_cond;
     t8_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue;
     t8_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output := t8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;

     -- n8_MUX[uxn_opcodes_h_l806_c7_1307] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l806_c7_1307_cond <= VAR_n8_MUX_uxn_opcodes_h_l806_c7_1307_cond;
     n8_MUX_uxn_opcodes_h_l806_c7_1307_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l806_c7_1307_iftrue;
     n8_MUX_uxn_opcodes_h_l806_c7_1307_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l806_c7_1307_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l806_c7_1307_return_output := n8_MUX_uxn_opcodes_h_l806_c7_1307_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l806_c7_1307] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l809_c7_0507] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse := VAR_n8_MUX_uxn_opcodes_h_l806_c7_1307_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l809_c7_0507_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l809_c7_0507_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l809_c7_0507_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l806_c7_1307_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l806_c7_1307_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l798_c2_0643_iffalse := VAR_t8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l803_c7_90ad] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l803_c7_90ad] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l806_c7_1307] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_return_output;

     -- t8_MUX[uxn_opcodes_h_l798_c2_0643] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l798_c2_0643_cond <= VAR_t8_MUX_uxn_opcodes_h_l798_c2_0643_cond;
     t8_MUX_uxn_opcodes_h_l798_c2_0643_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l798_c2_0643_iftrue;
     t8_MUX_uxn_opcodes_h_l798_c2_0643_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l798_c2_0643_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l798_c2_0643_return_output := t8_MUX_uxn_opcodes_h_l798_c2_0643_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l803_c7_90ad] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_cond;
     result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_return_output := result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l806_c7_1307] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_return_output;

     -- n8_MUX[uxn_opcodes_h_l803_c7_90ad] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l803_c7_90ad_cond <= VAR_n8_MUX_uxn_opcodes_h_l803_c7_90ad_cond;
     n8_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue;
     n8_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output := n8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l806_c7_1307] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l798_c2_0643_iffalse := VAR_n8_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l806_c7_1307_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l806_c7_1307_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l806_c7_1307_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l798_c2_0643_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l803_c7_90ad] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l798_c2_0643] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l798_c2_0643] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_cond;
     result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_return_output := result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l803_c7_90ad] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;

     -- n8_MUX[uxn_opcodes_h_l798_c2_0643] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l798_c2_0643_cond <= VAR_n8_MUX_uxn_opcodes_h_l798_c2_0643_cond;
     n8_MUX_uxn_opcodes_h_l798_c2_0643_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l798_c2_0643_iftrue;
     n8_MUX_uxn_opcodes_h_l798_c2_0643_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l798_c2_0643_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l798_c2_0643_return_output := n8_MUX_uxn_opcodes_h_l798_c2_0643_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l798_c2_0643] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l803_c7_90ad] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l798_c2_0643_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l803_c7_90ad_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l798_c2_0643] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l798_c2_0643] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l798_c2_0643] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l823_l794_DUPLICATE_89d4 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l823_l794_DUPLICATE_89d4_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l798_c2_0643_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l798_c2_0643_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l798_c2_0643_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l798_c2_0643_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l798_c2_0643_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l823_l794_DUPLICATE_89d4_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l823_l794_DUPLICATE_89d4_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
