-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity gth_0CLK_441a128d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end gth_0CLK_441a128d;
architecture arch of gth_0CLK_441a128d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1810_c6_a2e1]
signal BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1810_c2_810a]
signal n8_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1810_c2_810a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1810_c2_810a]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1810_c2_810a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1810_c2_810a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1810_c2_810a]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1810_c2_810a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1810_c2_810a]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1810_c2_810a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1810_c2_810a]
signal result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1810_c2_810a]
signal t8_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1823_c11_35b4]
signal BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1823_c7_cda4]
signal n8_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1823_c7_cda4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1823_c7_cda4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1823_c7_cda4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1823_c7_cda4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1823_c7_cda4]
signal result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1823_c7_cda4]
signal t8_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1826_c11_96c9]
signal BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1826_c7_e007]
signal n8_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1826_c7_e007]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1826_c7_e007]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1826_c7_e007]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1826_c7_e007]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1826_c7_e007]
signal result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1826_c7_e007]
signal t8_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1829_c11_8cba]
signal BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1829_c7_eaed]
signal n8_MUX_uxn_opcodes_h_l1829_c7_eaed_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1829_c7_eaed]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1829_c7_eaed]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1829_c7_eaed]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1829_c7_eaed]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1829_c7_eaed]
signal result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1831_c30_f1b3]
signal sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_return_output : signed(3 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1834_c21_4a39]
signal BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_right : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1834_c21_9341]
signal MUX_uxn_opcodes_h_l1834_c21_9341_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1834_c21_9341_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1834_c21_9341_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1834_c21_9341_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_04b4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1
BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_left,
BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_right,
BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output);

-- n8_MUX_uxn_opcodes_h_l1810_c2_810a
n8_MUX_uxn_opcodes_h_l1810_c2_810a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1810_c2_810a_cond,
n8_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue,
n8_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse,
n8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a
result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a
result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a
result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a
result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a
result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a
result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_return_output);

-- t8_MUX_uxn_opcodes_h_l1810_c2_810a
t8_MUX_uxn_opcodes_h_l1810_c2_810a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1810_c2_810a_cond,
t8_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue,
t8_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse,
t8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4
BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_left,
BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_right,
BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_return_output);

-- n8_MUX_uxn_opcodes_h_l1823_c7_cda4
n8_MUX_uxn_opcodes_h_l1823_c7_cda4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1823_c7_cda4_cond,
n8_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue,
n8_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse,
n8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4
result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4
result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4
result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output);

-- t8_MUX_uxn_opcodes_h_l1823_c7_cda4
t8_MUX_uxn_opcodes_h_l1823_c7_cda4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1823_c7_cda4_cond,
t8_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue,
t8_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse,
t8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9
BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_left,
BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_right,
BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_return_output);

-- n8_MUX_uxn_opcodes_h_l1826_c7_e007
n8_MUX_uxn_opcodes_h_l1826_c7_e007 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1826_c7_e007_cond,
n8_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue,
n8_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse,
n8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007
result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_cond,
result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_return_output);

-- t8_MUX_uxn_opcodes_h_l1826_c7_e007
t8_MUX_uxn_opcodes_h_l1826_c7_e007 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1826_c7_e007_cond,
t8_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue,
t8_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse,
t8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba
BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_left,
BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_right,
BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_return_output);

-- n8_MUX_uxn_opcodes_h_l1829_c7_eaed
n8_MUX_uxn_opcodes_h_l1829_c7_eaed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1829_c7_eaed_cond,
n8_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue,
n8_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse,
n8_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed
result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed
result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed
result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed
result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_cond,
result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3
sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_ins,
sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_x,
sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_y,
sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39
BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39 : entity work.BIN_OP_GT_uint8_t_uint8_t_0CLK_380ecc95 port map (
BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_left,
BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_right,
BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_return_output);

-- MUX_uxn_opcodes_h_l1834_c21_9341
MUX_uxn_opcodes_h_l1834_c21_9341 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1834_c21_9341_cond,
MUX_uxn_opcodes_h_l1834_c21_9341_iftrue,
MUX_uxn_opcodes_h_l1834_c21_9341_iffalse,
MUX_uxn_opcodes_h_l1834_c21_9341_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output,
 n8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
 t8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_return_output,
 n8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output,
 t8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_return_output,
 n8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_return_output,
 t8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_return_output,
 n8_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output,
 sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_return_output,
 MUX_uxn_opcodes_h_l1834_c21_9341_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1820_c3_e6cb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1815_c3_9332 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1810_c2_810a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1824_c3_5aae : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1823_c7_cda4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1826_c7_e007_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1829_c7_eaed_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1833_c3_dafb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1834_c21_9341_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1834_c21_9341_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1834_c21_9341_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1834_c21_9341_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1823_l1826_l1810_l1829_DUPLICATE_7608_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_1255_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_8613_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_ec16_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1826_l1829_DUPLICATE_254a_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1838_l1806_DUPLICATE_bcb3_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1833_c3_dafb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1833_c3_dafb;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1824_c3_5aae := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1824_c3_5aae;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1834_c21_9341_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1815_c3_9332 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1815_c3_9332;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_right := to_unsigned(2, 2);
     VAR_MUX_uxn_opcodes_h_l1834_c21_9341_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1820_c3_e6cb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1820_c3_e6cb;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse := t8;
     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1810_c2_810a_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_1255 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_1255_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1823_l1826_l1810_l1829_DUPLICATE_7608 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1823_l1826_l1810_l1829_DUPLICATE_7608_return_output := result.u8_value;

     -- BIN_OP_GT[uxn_opcodes_h_l1834_c21_4a39] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_left;
     BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_return_output := BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1826_c11_96c9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_ec16 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_ec16_return_output := result.is_stack_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1810_c2_810a_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1829_c11_8cba] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_left;
     BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_return_output := BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1826_l1829_DUPLICATE_254a LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1826_l1829_DUPLICATE_254a_return_output := result.stack_address_sp_offset;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1810_c2_810a_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_8613 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_8613_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l1831_c30_f1b3] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_ins;
     sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_x;
     sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_return_output := sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1810_c2_810a_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1810_c6_a2e1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1823_c11_35b4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1810_c2_810a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1810_c2_810a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1810_c6_a2e1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1823_c7_cda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1823_c7_cda4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1823_c11_35b4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1826_c7_e007_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1826_c7_e007_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c11_96c9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1829_c7_eaed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1829_c11_8cba_return_output;
     VAR_MUX_uxn_opcodes_h_l1834_c21_9341_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1834_c21_4a39_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_1255_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_1255_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_1255_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_8613_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_8613_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_8613_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_ec16_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_ec16_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1823_l1826_l1829_DUPLICATE_ec16_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1826_l1829_DUPLICATE_254a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1826_l1829_DUPLICATE_254a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1823_l1826_l1810_l1829_DUPLICATE_7608_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1823_l1826_l1810_l1829_DUPLICATE_7608_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1823_l1826_l1810_l1829_DUPLICATE_7608_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1823_l1826_l1810_l1829_DUPLICATE_7608_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1810_c2_810a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1810_c2_810a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1810_c2_810a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1810_c2_810a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1831_c30_f1b3_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1829_c7_eaed] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output;

     -- n8_MUX[uxn_opcodes_h_l1829_c7_eaed] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1829_c7_eaed_cond <= VAR_n8_MUX_uxn_opcodes_h_l1829_c7_eaed_cond;
     n8_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue;
     n8_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output := n8_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1829_c7_eaed] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1829_c7_eaed] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output;

     -- MUX[uxn_opcodes_h_l1834_c21_9341] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1834_c21_9341_cond <= VAR_MUX_uxn_opcodes_h_l1834_c21_9341_cond;
     MUX_uxn_opcodes_h_l1834_c21_9341_iftrue <= VAR_MUX_uxn_opcodes_h_l1834_c21_9341_iftrue;
     MUX_uxn_opcodes_h_l1834_c21_9341_iffalse <= VAR_MUX_uxn_opcodes_h_l1834_c21_9341_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1834_c21_9341_return_output := MUX_uxn_opcodes_h_l1834_c21_9341_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1829_c7_eaed] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_return_output;

     -- t8_MUX[uxn_opcodes_h_l1826_c7_e007] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1826_c7_e007_cond <= VAR_t8_MUX_uxn_opcodes_h_l1826_c7_e007_cond;
     t8_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue;
     t8_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output := t8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue := VAR_MUX_uxn_opcodes_h_l1834_c21_9341_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;
     -- n8_MUX[uxn_opcodes_h_l1826_c7_e007] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1826_c7_e007_cond <= VAR_n8_MUX_uxn_opcodes_h_l1826_c7_e007_cond;
     n8_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue;
     n8_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output := n8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1826_c7_e007] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;

     -- t8_MUX[uxn_opcodes_h_l1823_c7_cda4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1823_c7_cda4_cond <= VAR_t8_MUX_uxn_opcodes_h_l1823_c7_cda4_cond;
     t8_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue;
     t8_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output := t8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1826_c7_e007] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1826_c7_e007] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1829_c7_eaed] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output := result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1826_c7_e007] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1829_c7_eaed_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1823_c7_cda4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1823_c7_cda4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1826_c7_e007] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_return_output := result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;

     -- t8_MUX[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1810_c2_810a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1810_c2_810a_cond;
     t8_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue;
     t8_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output := t8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1823_c7_cda4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1823_c7_cda4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1823_c7_cda4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1823_c7_cda4_cond <= VAR_n8_MUX_uxn_opcodes_h_l1823_c7_cda4_cond;
     n8_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue;
     n8_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output := n8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c7_e007_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output;

     -- n8_MUX[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1810_c2_810a_cond <= VAR_n8_MUX_uxn_opcodes_h_l1810_c2_810a_cond;
     n8_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue;
     n8_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output := n8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1823_c7_cda4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1810_c2_810a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1823_c7_cda4_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1810_c2_810a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1838_l1806_DUPLICATE_bcb3 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1838_l1806_DUPLICATE_bcb3_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_04b4(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1810_c2_810a_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1810_c2_810a_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1838_l1806_DUPLICATE_bcb3_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1838_l1806_DUPLICATE_bcb3_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
