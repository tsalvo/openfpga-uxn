-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 37
entity dup_0CLK_6be78140 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_6be78140;
architecture arch of dup_0CLK_6be78140 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2620_c6_a200]
signal BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2620_c1_dcb5]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2620_c2_240d]
signal t8_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2620_c2_240d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2620_c2_240d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2620_c2_240d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2620_c2_240d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2620_c2_240d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2620_c2_240d]
signal result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2621_c3_d2d5[uxn_opcodes_h_l2621_c3_d2d5]
signal printf_uxn_opcodes_h_l2621_c3_d2d5_uxn_opcodes_h_l2621_c3_d2d5_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2625_c11_b631]
signal BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2625_c7_3417]
signal t8_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2625_c7_3417]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2625_c7_3417]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2625_c7_3417]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2625_c7_3417]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2625_c7_3417]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2625_c7_3417]
signal result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2628_c11_a19a]
signal BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2628_c7_b5b2]
signal t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2628_c7_b5b2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2628_c7_b5b2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2628_c7_b5b2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2628_c7_b5b2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2628_c7_b5b2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2628_c7_b5b2]
signal result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2631_c30_69e1]
signal sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2636_c11_8d7c]
signal BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2636_c7_ff17]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2636_c7_ff17]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2636_c7_ff17]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2636_c7_ff17]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2636_c7_ff17]
signal result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2641_c11_371a]
signal BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2641_c7_c2b8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2641_c7_c2b8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_4e73( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200
BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_left,
BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_right,
BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_return_output);

-- t8_MUX_uxn_opcodes_h_l2620_c2_240d
t8_MUX_uxn_opcodes_h_l2620_c2_240d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2620_c2_240d_cond,
t8_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue,
t8_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse,
t8_MUX_uxn_opcodes_h_l2620_c2_240d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d
result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d
result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_return_output);

-- printf_uxn_opcodes_h_l2621_c3_d2d5_uxn_opcodes_h_l2621_c3_d2d5
printf_uxn_opcodes_h_l2621_c3_d2d5_uxn_opcodes_h_l2621_c3_d2d5 : entity work.printf_uxn_opcodes_h_l2621_c3_d2d5_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2621_c3_d2d5_uxn_opcodes_h_l2621_c3_d2d5_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631
BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_left,
BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_right,
BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_return_output);

-- t8_MUX_uxn_opcodes_h_l2625_c7_3417
t8_MUX_uxn_opcodes_h_l2625_c7_3417 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2625_c7_3417_cond,
t8_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue,
t8_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse,
t8_MUX_uxn_opcodes_h_l2625_c7_3417_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417
result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417
result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417
result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417
result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417
result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_cond,
result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a
BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_left,
BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_right,
BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_return_output);

-- t8_MUX_uxn_opcodes_h_l2628_c7_b5b2
t8_MUX_uxn_opcodes_h_l2628_c7_b5b2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond,
t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue,
t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse,
t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2
result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2
result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2
result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2
result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1
sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_ins,
sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_x,
sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_y,
sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c
BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_left,
BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_right,
BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17
result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17
result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17
result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17
result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_cond,
result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a
BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_left,
BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_right,
BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8
result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8
result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_return_output,
 t8_MUX_uxn_opcodes_h_l2620_c2_240d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_return_output,
 t8_MUX_uxn_opcodes_h_l2625_c7_3417_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_return_output,
 t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output,
 sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2622_c3_46a0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2621_c3_d2d5_uxn_opcodes_h_l2621_c3_d2d5_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2626_c3_0eaa : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2633_c3_9a13 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2638_c3_ae29 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2636_c7_ff17_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2620_l2636_l2625_l2641_DUPLICATE_8727_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2620_l2636_l2625_DUPLICATE_5ed4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2620_l2625_l2628_DUPLICATE_4afb_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2620_l2636_l2625_DUPLICATE_447b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2636_l2625_l2641_l2628_DUPLICATE_9988_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l2646_l2616_DUPLICATE_0822_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2622_c3_46a0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2622_c3_46a0;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2633_c3_9a13 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2633_c3_9a13;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2626_c3_0eaa := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2626_c3_0eaa;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2638_c3_ae29 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2638_c3_ae29;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_iffalse := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l2631_c30_69e1] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_ins;
     sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_x;
     sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_return_output := sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2628_c11_a19a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2620_l2625_l2628_DUPLICATE_4afb LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2620_l2625_l2628_DUPLICATE_4afb_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2641_c11_371a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2636_c11_8d7c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2625_c11_b631] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_left;
     BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_return_output := BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2620_l2636_l2625_DUPLICATE_447b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2620_l2636_l2625_DUPLICATE_447b_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2620_l2636_l2625_DUPLICATE_5ed4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2620_l2636_l2625_DUPLICATE_5ed4_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2620_c6_a200] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_left;
     BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output := BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2620_l2636_l2625_l2641_DUPLICATE_8727 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2620_l2636_l2625_l2641_DUPLICATE_8727_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2636_l2625_l2641_l2628_DUPLICATE_9988 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2636_l2625_l2641_l2628_DUPLICATE_9988_return_output := result.is_opc_done;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2636_c7_ff17] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2636_c7_ff17_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2620_c2_240d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2620_c6_a200_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2625_c7_3417_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2625_c11_b631_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2628_c11_a19a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2636_c11_8d7c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2641_c11_371a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2620_l2625_l2628_DUPLICATE_4afb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2620_l2625_l2628_DUPLICATE_4afb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2620_l2625_l2628_DUPLICATE_4afb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2636_l2625_l2641_l2628_DUPLICATE_9988_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2636_l2625_l2641_l2628_DUPLICATE_9988_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2636_l2625_l2641_l2628_DUPLICATE_9988_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2636_l2625_l2641_l2628_DUPLICATE_9988_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2620_l2636_l2625_DUPLICATE_5ed4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2620_l2636_l2625_DUPLICATE_5ed4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2620_l2636_l2625_DUPLICATE_5ed4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2620_l2636_l2625_l2641_DUPLICATE_8727_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2620_l2636_l2625_l2641_DUPLICATE_8727_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2620_l2636_l2625_l2641_DUPLICATE_8727_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2620_l2636_l2625_l2641_DUPLICATE_8727_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2620_l2636_l2625_DUPLICATE_447b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2620_l2636_l2625_DUPLICATE_447b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2620_l2636_l2625_DUPLICATE_447b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2636_c7_ff17_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2631_c30_69e1_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2628_c7_b5b2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2620_c1_dcb5] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2636_c7_ff17] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2641_c7_c2b8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2636_c7_ff17] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output;

     -- t8_MUX[uxn_opcodes_h_l2628_c7_b5b2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond <= VAR_t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond;
     t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue;
     t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output := t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2641_c7_c2b8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2636_c7_ff17] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output := result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2621_c3_d2d5_uxn_opcodes_h_l2621_c3_d2d5_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2620_c1_dcb5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2641_c7_c2b8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;
     -- t8_MUX[uxn_opcodes_h_l2625_c7_3417] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2625_c7_3417_cond <= VAR_t8_MUX_uxn_opcodes_h_l2625_c7_3417_cond;
     t8_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue;
     t8_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2625_c7_3417_return_output := t8_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2628_c7_b5b2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2625_c7_3417] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2636_c7_ff17] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2628_c7_b5b2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;

     -- printf_uxn_opcodes_h_l2621_c3_d2d5[uxn_opcodes_h_l2621_c3_d2d5] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2621_c3_d2d5_uxn_opcodes_h_l2621_c3_d2d5_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2621_c3_d2d5_uxn_opcodes_h_l2621_c3_d2d5_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2628_c7_b5b2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2636_c7_ff17] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2636_c7_ff17_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2625_c7_3417] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2625_c7_3417] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2628_c7_b5b2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2625_c7_3417] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_return_output := result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2628_c7_b5b2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;

     -- t8_MUX[uxn_opcodes_h_l2620_c2_240d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2620_c2_240d_cond <= VAR_t8_MUX_uxn_opcodes_h_l2620_c2_240d_cond;
     t8_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue;
     t8_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2620_c2_240d_return_output := t8_MUX_uxn_opcodes_h_l2620_c2_240d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2620_c2_240d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2628_c7_b5b2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2620_c2_240d_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2625_c7_3417] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2620_c2_240d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2625_c7_3417] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2620_c2_240d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2620_c2_240d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2625_c7_3417_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2620_c2_240d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2620_c2_240d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l2646_l2616_DUPLICATE_0822 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l2646_l2616_DUPLICATE_0822_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4e73(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2620_c2_240d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2620_c2_240d_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2620_c2_240d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2620_c2_240d_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2620_c2_240d_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l2646_l2616_DUPLICATE_0822_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l2646_l2616_DUPLICATE_0822_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
