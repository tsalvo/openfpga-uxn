-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 114
entity deo2_0CLK_0f83c89f is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_device_ram_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end deo2_0CLK_0f83c89f;
architecture arch of deo2_0CLK_0f83c89f is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal current_deo_phase : unsigned(7 downto 0) := to_unsigned(0, 8);
signal deo_param0 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal deo_param1 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal is_second_deo : unsigned(0 downto 0) := to_unsigned(0, 1);
signal result : opcode_result_t := opcode_result_t_NULL;
signal device_out_result : device_out_result_t := device_out_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_current_deo_phase : unsigned(7 downto 0);
signal REG_COMB_deo_param0 : unsigned(7 downto 0);
signal REG_COMB_deo_param1 : unsigned(7 downto 0);
signal REG_COMB_is_second_deo : unsigned(0 downto 0);
signal REG_COMB_result : opcode_result_t;
signal REG_COMB_device_out_result : device_out_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l533_c6_ea52]
signal BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l533_c1_1764]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);

-- deo_param1_MUX[uxn_opcodes_h_l533_c2_51df]
signal deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l533_c2_51df]
signal l8_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l533_c2_51df]
signal t8_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l533_c2_51df]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l533_c2_51df]
signal result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(15 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l533_c2_51df]
signal result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l533_c2_51df]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(3 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l533_c2_51df]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(0 downto 0);

-- result_vram_address_MUX[uxn_opcodes_h_l533_c2_51df]
signal result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(31 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(31 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(31 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l533_c2_51df]
signal result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l533_c2_51df]
signal result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l533_c2_51df]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l533_c2_51df]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l533_c2_51df]
signal result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l533_c2_51df]
signal n8_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l533_c2_51df]
signal device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_return_output : device_out_result_t;

-- deo_param0_MUX[uxn_opcodes_h_l533_c2_51df]
signal deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l533_c2_51df]
signal current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l533_c2_51df]
signal is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l534_c3_7035[uxn_opcodes_h_l534_c3_7035]
signal printf_uxn_opcodes_h_l534_c3_7035_uxn_opcodes_h_l534_c3_7035_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l540_c11_f922]
signal BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l543_c7_d631]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);

-- deo_param1_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal l8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal t8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(15 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(3 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);

-- result_vram_address_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(31 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(31 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(31 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal n8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : device_out_result_t;

-- deo_param0_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l540_c7_7e3c]
signal is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l543_c11_61df]
signal BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);

-- deo_param1_MUX[uxn_opcodes_h_l543_c7_d631]
signal deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l543_c7_d631]
signal l8_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l543_c7_d631]
signal t8_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l543_c7_d631]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l543_c7_d631]
signal result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(15 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l543_c7_d631]
signal result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l543_c7_d631]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(3 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l543_c7_d631]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);

-- result_vram_address_MUX[uxn_opcodes_h_l543_c7_d631]
signal result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(31 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(31 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(31 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l543_c7_d631]
signal result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l543_c7_d631]
signal result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l543_c7_d631]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l543_c7_d631]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l543_c7_d631]
signal result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l543_c7_d631]
signal n8_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l543_c7_d631]
signal device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_return_output : device_out_result_t;

-- deo_param0_MUX[uxn_opcodes_h_l543_c7_d631]
signal deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l543_c7_d631]
signal current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l543_c7_d631]
signal is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l547_c11_ed5d]
signal BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l550_c7_c749]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);

-- deo_param1_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal l8_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(15 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(3 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);

-- result_vram_address_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(31 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(31 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(31 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal n8_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : device_out_result_t;

-- deo_param0_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l547_c7_f1ac]
signal is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l550_c11_a93d]
signal BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l556_c1_7044]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_return_output : unsigned(0 downto 0);

-- deo_param1_MUX[uxn_opcodes_h_l550_c7_c749]
signal deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l550_c7_c749]
signal l8_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l550_c7_c749]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l550_c7_c749]
signal result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(15 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l550_c7_c749]
signal result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l550_c7_c749]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(3 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l550_c7_c749]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);

-- result_vram_address_MUX[uxn_opcodes_h_l550_c7_c749]
signal result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(31 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(31 downto 0);
signal result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(31 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l550_c7_c749]
signal result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l550_c7_c749]
signal result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l550_c7_c749]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l550_c7_c749]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l550_c7_c749]
signal result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(7 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l550_c7_c749]
signal device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_return_output : device_out_result_t;

-- deo_param0_MUX[uxn_opcodes_h_l550_c7_c749]
signal deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(7 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l550_c7_c749]
signal current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(7 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l550_c7_c749]
signal is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l554_c30_0d04]
signal sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l558_c32_4775]
signal BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_return_output : unsigned(8 downto 0);

-- MUX[uxn_opcodes_h_l558_c16_1f6e]
signal MUX_uxn_opcodes_h_l558_c16_1f6e_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l558_c16_1f6e_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l558_c16_1f6e_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l558_c16_1f6e_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l559_c16_91f7]
signal MUX_uxn_opcodes_h_l559_c16_91f7_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l559_c16_91f7_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l559_c16_91f7_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l559_c16_91f7_return_output : unsigned(7 downto 0);

-- device_out[uxn_opcodes_h_l560_c23_82e8]
signal device_out_uxn_opcodes_h_l560_c23_82e8_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_out_uxn_opcodes_h_l560_c23_82e8_device_address : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l560_c23_82e8_value : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l560_c23_82e8_phase : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l560_c23_82e8_previous_device_ram_read : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l560_c23_82e8_previous_ram_read : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l560_c23_82e8_return_output : device_out_result_t;

-- BIN_OP_AND[uxn_opcodes_h_l568_c24_9a70]
signal BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_left : unsigned(0 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_right : unsigned(0 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_return_output : unsigned(0 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l569_c3_57f7]
signal current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_return_output : unsigned(7 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l569_c3_57f7]
signal is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l573_c4_0b8c]
signal BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_return_output : unsigned(8 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e309( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : signed;
 ref_toks_11 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_sp_shift := ref_toks_1;
      base.u16_value := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.vram_write_layer := ref_toks_5;
      base.vram_address := ref_toks_6;
      base.device_ram_address := ref_toks_7;
      base.is_opc_done := ref_toks_8;
      base.is_device_ram_write := ref_toks_9;
      base.sp_relative_shift := ref_toks_10;
      base.u8_value := ref_toks_11;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52
BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_left,
BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_right,
BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- deo_param1_MUX_uxn_opcodes_h_l533_c2_51df
deo_param1_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_cond,
deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- l8_MUX_uxn_opcodes_h_l533_c2_51df
l8_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l533_c2_51df_cond,
l8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
l8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
l8_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- t8_MUX_uxn_opcodes_h_l533_c2_51df
t8_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l533_c2_51df_cond,
t8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
t8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
t8_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df
result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df
result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_cond,
result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df
result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df
result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df
result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_cond,
result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df
result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df
result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df
result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df
result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df
result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_cond,
result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- n8_MUX_uxn_opcodes_h_l533_c2_51df
n8_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l533_c2_51df_cond,
n8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
n8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
n8_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l533_c2_51df
device_out_result_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_cond,
device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- deo_param0_MUX_uxn_opcodes_h_l533_c2_51df
deo_param0_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_cond,
deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df
current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_cond,
current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df
is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_cond,
is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

-- printf_uxn_opcodes_h_l534_c3_7035_uxn_opcodes_h_l534_c3_7035
printf_uxn_opcodes_h_l534_c3_7035_uxn_opcodes_h_l534_c3_7035 : entity work.printf_uxn_opcodes_h_l534_c3_7035_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l534_c3_7035_uxn_opcodes_h_l534_c3_7035_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922
BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_left,
BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_right,
BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c
deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- l8_MUX_uxn_opcodes_h_l540_c7_7e3c
l8_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
l8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
l8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
l8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- t8_MUX_uxn_opcodes_h_l540_c7_7e3c
t8_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
t8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
t8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
t8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c
result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c
result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c
result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c
result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c
result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c
result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c
result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c
result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c
result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c
result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- n8_MUX_uxn_opcodes_h_l540_c7_7e3c
n8_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
n8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
n8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
n8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c
device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c
deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c
current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c
is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_cond,
is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df
BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_left,
BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_right,
BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- deo_param1_MUX_uxn_opcodes_h_l543_c7_d631
deo_param1_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_cond,
deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- l8_MUX_uxn_opcodes_h_l543_c7_d631
l8_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l543_c7_d631_cond,
l8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
l8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
l8_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- t8_MUX_uxn_opcodes_h_l543_c7_d631
t8_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l543_c7_d631_cond,
t8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
t8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
t8_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631
result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631
result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_cond,
result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631
result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631
result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631
result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_cond,
result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631
result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631
result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631
result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631
result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631
result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_cond,
result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- n8_MUX_uxn_opcodes_h_l543_c7_d631
n8_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l543_c7_d631_cond,
n8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
n8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
n8_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l543_c7_d631
device_out_result_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_cond,
device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- deo_param0_MUX_uxn_opcodes_h_l543_c7_d631
deo_param0_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_cond,
deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631
current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_cond,
current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631
is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_cond,
is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d
BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_left,
BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_right,
BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac
deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- l8_MUX_uxn_opcodes_h_l547_c7_f1ac
l8_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
l8_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
l8_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
l8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac
result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac
result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac
result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac
result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac
result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac
result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac
result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac
result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac
result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac
result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- n8_MUX_uxn_opcodes_h_l547_c7_f1ac
n8_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
n8_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
n8_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
n8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac
device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac
deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac
current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac
is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_cond,
is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d
BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_left,
BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_right,
BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_return_output);

-- deo_param1_MUX_uxn_opcodes_h_l550_c7_c749
deo_param1_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_cond,
deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- l8_MUX_uxn_opcodes_h_l550_c7_c749
l8_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l550_c7_c749_cond,
l8_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
l8_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
l8_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749
result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749
result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_cond,
result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749
result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749
result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749
result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_cond,
result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749
result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749
result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749
result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749
result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749
result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_cond,
result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l550_c7_c749
device_out_result_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_cond,
device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- deo_param0_MUX_uxn_opcodes_h_l550_c7_c749
deo_param0_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_cond,
deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749
current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_cond,
current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749
is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_cond,
is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_return_output);

-- sp_relative_shift_uxn_opcodes_h_l554_c30_0d04
sp_relative_shift_uxn_opcodes_h_l554_c30_0d04 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_ins,
sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_x,
sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_y,
sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775
BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_left,
BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_right,
BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_return_output);

-- MUX_uxn_opcodes_h_l558_c16_1f6e
MUX_uxn_opcodes_h_l558_c16_1f6e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l558_c16_1f6e_cond,
MUX_uxn_opcodes_h_l558_c16_1f6e_iftrue,
MUX_uxn_opcodes_h_l558_c16_1f6e_iffalse,
MUX_uxn_opcodes_h_l558_c16_1f6e_return_output);

-- MUX_uxn_opcodes_h_l559_c16_91f7
MUX_uxn_opcodes_h_l559_c16_91f7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l559_c16_91f7_cond,
MUX_uxn_opcodes_h_l559_c16_91f7_iftrue,
MUX_uxn_opcodes_h_l559_c16_91f7_iffalse,
MUX_uxn_opcodes_h_l559_c16_91f7_return_output);

-- device_out_uxn_opcodes_h_l560_c23_82e8
device_out_uxn_opcodes_h_l560_c23_82e8 : entity work.device_out_0CLK_f5486376 port map (
clk,
device_out_uxn_opcodes_h_l560_c23_82e8_CLOCK_ENABLE,
device_out_uxn_opcodes_h_l560_c23_82e8_device_address,
device_out_uxn_opcodes_h_l560_c23_82e8_value,
device_out_uxn_opcodes_h_l560_c23_82e8_phase,
device_out_uxn_opcodes_h_l560_c23_82e8_previous_device_ram_read,
device_out_uxn_opcodes_h_l560_c23_82e8_previous_ram_read,
device_out_uxn_opcodes_h_l560_c23_82e8_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70
BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_left,
BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_right,
BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7
current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_cond,
current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7
is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_cond,
is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c
BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_left,
BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_right,
BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_device_ram_read,
 previous_ram_read,
 -- Registers
 t8,
 n8,
 l8,
 current_deo_phase,
 deo_param0,
 deo_param1,
 is_second_deo,
 result,
 device_out_result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 l8_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 t8_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 n8_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 l8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 t8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 n8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 l8_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 t8_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 n8_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 l8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 n8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_return_output,
 deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 l8_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_return_output,
 sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_return_output,
 MUX_uxn_opcodes_h_l558_c16_1f6e_return_output,
 MUX_uxn_opcodes_h_l559_c16_91f7_return_output,
 device_out_uxn_opcodes_h_l560_c23_82e8_return_output,
 BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l535_c3_25fe : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_uxn_opcodes_h_l538_c3_92e4 : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l534_c3_7035_uxn_opcodes_h_l534_c3_7035_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l541_c3_c98c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l544_c3_32b3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_iffalse : unsigned(0 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l552_c3_01c0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(31 downto 0);
 variable VAR_result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l558_c16_1f6e_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l558_c16_1f6e_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l558_c16_1f6e_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_return_output : unsigned(8 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l558_c16_1f6e_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l559_c16_91f7_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l559_c16_91f7_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l559_c16_91f7_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l559_c16_91f7_return_output : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l560_c23_82e8_device_address : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l560_c23_82e8_value : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l560_c23_82e8_phase : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l560_c23_82e8_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l560_c23_82e8_previous_ram_read : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l560_c23_82e8_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l560_c23_82e8_return_output : device_out_result_t;
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l561_c32_e0b2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l562_c31_8d15_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l563_c26_a98f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l564_c29_faf0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_device_out_result_t_vram_address_d41d_uxn_opcodes_h_l565_c25_61d4_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_device_out_result_t_ram_address_d41d_uxn_opcodes_h_l566_c22_dca3_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l567_c21_c2b2_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_return_output : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_uxn_opcodes_h_l570_c4_3f4b : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_uxn_opcodes_h_l573_c4_bcfc : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_cond : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_return_output : unsigned(8 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l543_l533_l547_l540_DUPLICATE_f70a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_2129_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_5740_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b34b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_opcode_result_t_vram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_11c0_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b4bc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_cf78_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_aa12_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_d12a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l543_l547_l540_l550_DUPLICATE_0003_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l547_l550_DUPLICATE_8042_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l568_l569_DUPLICATE_6038_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e309_uxn_opcodes_h_l577_l527_DUPLICATE_9675_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_current_deo_phase : unsigned(7 downto 0);
variable REG_VAR_deo_param0 : unsigned(7 downto 0);
variable REG_VAR_deo_param1 : unsigned(7 downto 0);
variable REG_VAR_is_second_deo : unsigned(0 downto 0);
variable REG_VAR_result : opcode_result_t;
variable REG_VAR_device_out_result : device_out_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_current_deo_phase := current_deo_phase;
  REG_VAR_deo_param0 := deo_param0;
  REG_VAR_deo_param1 := deo_param1;
  REG_VAR_is_second_deo := is_second_deo;
  REG_VAR_result := result;
  REG_VAR_device_out_result := device_out_result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_right := to_unsigned(2, 2);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_right := to_unsigned(0, 1);
     VAR_is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_current_deo_phase_uxn_opcodes_h_l538_c3_92e4 := resize(to_unsigned(0, 1), 8);
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := VAR_current_deo_phase_uxn_opcodes_h_l538_c3_92e4;
     VAR_current_deo_phase_uxn_opcodes_h_l570_c4_3f4b := resize(to_unsigned(0, 1), 8);
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_iftrue := VAR_current_deo_phase_uxn_opcodes_h_l570_c4_3f4b;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l535_c3_25fe := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l535_c3_25fe;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := to_unsigned(0, 1);
     VAR_is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_y := resize(to_signed(-3, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l541_c3_c98c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l541_c3_c98c;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l544_c3_32b3 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l544_c3_32b3;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l552_c3_01c0 := resize(to_unsigned(0, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l552_c3_01c0;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_device_ram_read := previous_device_ram_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_left := current_deo_phase;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := current_deo_phase;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := current_deo_phase;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := current_deo_phase;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := current_deo_phase;
     VAR_device_out_uxn_opcodes_h_l560_c23_82e8_phase := current_deo_phase;
     VAR_deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := deo_param0;
     VAR_deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := deo_param0;
     VAR_deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := deo_param0;
     VAR_deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := deo_param0;
     VAR_deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := deo_param0;
     VAR_deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := deo_param1;
     VAR_deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := deo_param1;
     VAR_deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := deo_param1;
     VAR_deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := deo_param1;
     VAR_deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := deo_param1;
     VAR_device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := device_out_result;
     VAR_device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := device_out_result;
     VAR_device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := device_out_result;
     VAR_device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := device_out_result;
     VAR_device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := device_out_result;
     VAR_sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_ins := VAR_ins;
     VAR_BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_right := is_second_deo;
     VAR_MUX_uxn_opcodes_h_l558_c16_1f6e_cond := is_second_deo;
     VAR_MUX_uxn_opcodes_h_l559_c16_91f7_cond := is_second_deo;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := is_second_deo;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := is_second_deo;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := is_second_deo;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := is_second_deo;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_iffalse := is_second_deo;
     VAR_MUX_uxn_opcodes_h_l559_c16_91f7_iffalse := l8;
     VAR_l8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := l8;
     VAR_MUX_uxn_opcodes_h_l559_c16_91f7_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_left := VAR_phase;
     VAR_device_out_uxn_opcodes_h_l560_c23_82e8_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_device_out_uxn_opcodes_h_l560_c23_82e8_previous_ram_read := VAR_previous_ram_read;
     VAR_l8_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_left := t8;
     VAR_MUX_uxn_opcodes_h_l558_c16_1f6e_iffalse := t8;
     VAR_t8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := t8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l547_l550_DUPLICATE_8042 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l547_l550_DUPLICATE_8042_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint32_t_opcode_result_t_vram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_11c0 LATENCY=0
     VAR_CONST_REF_RD_uint32_t_opcode_result_t_vram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_11c0_return_output := result.vram_address;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_d12a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_d12a_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_cf78 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_cf78_return_output := result.is_device_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b34b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b34b_return_output := result.vram_write_layer;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l543_l547_l540_l550_DUPLICATE_0003 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l543_l547_l540_l550_DUPLICATE_0003_return_output := result.is_opc_done;

     -- BIN_OP_PLUS[uxn_opcodes_h_l558_c32_4775] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_left;
     BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_return_output := BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b4bc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b4bc_return_output := result.device_ram_address;

     -- BIN_OP_EQ[uxn_opcodes_h_l543_c11_61df] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_left;
     BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output := BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l554_c30_0d04] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_ins;
     sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_x <= VAR_sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_x;
     sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_y <= VAR_sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_return_output := sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l540_c11_f922] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_left;
     BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output := BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l547_c11_ed5d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_left;
     BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output := BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l533_c6_ea52] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_left;
     BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output := BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l573_c4_0b8c] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_left;
     BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_return_output := BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_aa12 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_aa12_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_5740 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_5740_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_2129 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_2129_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l550_c11_a93d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_left;
     BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output := BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l543_l533_l547_l540_DUPLICATE_f70a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l543_l533_l547_l540_DUPLICATE_f70a_return_output := result.is_sp_shift;

     -- MUX[uxn_opcodes_h_l559_c16_91f7] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l559_c16_91f7_cond <= VAR_MUX_uxn_opcodes_h_l559_c16_91f7_cond;
     MUX_uxn_opcodes_h_l559_c16_91f7_iftrue <= VAR_MUX_uxn_opcodes_h_l559_c16_91f7_iftrue;
     MUX_uxn_opcodes_h_l559_c16_91f7_iffalse <= VAR_MUX_uxn_opcodes_h_l559_c16_91f7_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l559_c16_91f7_return_output := MUX_uxn_opcodes_h_l559_c16_91f7_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l533_c2_51df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l533_c6_ea52_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l540_c11_f922_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l543_c7_d631_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l543_c11_61df_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l547_c11_ed5d_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l550_c11_a93d_return_output;
     VAR_MUX_uxn_opcodes_h_l558_c16_1f6e_iftrue := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l558_c32_4775_return_output, 8);
     VAR_current_deo_phase_uxn_opcodes_h_l573_c4_bcfc := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l573_c4_0b8c_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_aa12_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_aa12_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_aa12_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_aa12_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_aa12_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_2129_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_2129_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_2129_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_2129_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_2129_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_cf78_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_cf78_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_cf78_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_cf78_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_cf78_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l543_l547_l540_l550_DUPLICATE_0003_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l543_l547_l540_l550_DUPLICATE_0003_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l543_l547_l540_l550_DUPLICATE_0003_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l543_l547_l540_l550_DUPLICATE_0003_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l543_l533_l547_l540_DUPLICATE_f70a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l543_l533_l547_l540_DUPLICATE_f70a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l543_l533_l547_l540_DUPLICATE_f70a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l543_l533_l547_l540_DUPLICATE_f70a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_5740_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_5740_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_5740_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_5740_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_5740_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b34b_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b34b_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b34b_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b34b_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b34b_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := VAR_CONST_REF_RD_uint32_t_opcode_result_t_vram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_11c0_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := VAR_CONST_REF_RD_uint32_t_opcode_result_t_vram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_11c0_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := VAR_CONST_REF_RD_uint32_t_opcode_result_t_vram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_11c0_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := VAR_CONST_REF_RD_uint32_t_opcode_result_t_vram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_11c0_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := VAR_CONST_REF_RD_uint32_t_opcode_result_t_vram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_11c0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l547_l550_DUPLICATE_8042_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l547_l550_DUPLICATE_8042_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b4bc_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b4bc_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b4bc_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b4bc_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_b4bc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_d12a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_d12a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_d12a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_d12a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l550_l547_l543_l540_l533_DUPLICATE_d12a_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_MUX_uxn_opcodes_h_l559_c16_91f7_return_output;
     VAR_device_out_uxn_opcodes_h_l560_c23_82e8_value := VAR_MUX_uxn_opcodes_h_l559_c16_91f7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l554_c30_0d04_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_iffalse := VAR_current_deo_phase_uxn_opcodes_h_l573_c4_bcfc;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- deo_param1_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_return_output := deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- l8_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_l8_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     l8_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     l8_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l550_c7_c749_return_output := l8_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- n8_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_n8_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     n8_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     n8_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := n8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- MUX[uxn_opcodes_h_l558_c16_1f6e] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l558_c16_1f6e_cond <= VAR_MUX_uxn_opcodes_h_l558_c16_1f6e_cond;
     MUX_uxn_opcodes_h_l558_c16_1f6e_iftrue <= VAR_MUX_uxn_opcodes_h_l558_c16_1f6e_iftrue;
     MUX_uxn_opcodes_h_l558_c16_1f6e_iffalse <= VAR_MUX_uxn_opcodes_h_l558_c16_1f6e_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l558_c16_1f6e_return_output := MUX_uxn_opcodes_h_l558_c16_1f6e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- t8_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_t8_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     t8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     t8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l543_c7_d631_return_output := t8_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l533_c1_1764] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_MUX_uxn_opcodes_h_l558_c16_1f6e_return_output;
     VAR_device_out_uxn_opcodes_h_l560_c23_82e8_device_address := VAR_MUX_uxn_opcodes_h_l558_c16_1f6e_return_output;
     VAR_printf_uxn_opcodes_h_l534_c3_7035_uxn_opcodes_h_l534_c3_7035_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l533_c1_1764_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_deo_param1_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_l8_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_n8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     -- printf_uxn_opcodes_h_l534_c3_7035[uxn_opcodes_h_l534_c3_7035] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l534_c3_7035_uxn_opcodes_h_l534_c3_7035_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l534_c3_7035_uxn_opcodes_h_l534_c3_7035_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- n8_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_n8_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     n8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     n8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l543_c7_d631_return_output := n8_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- t8_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_t8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     t8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     t8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := t8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- deo_param0_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_return_output := deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- l8_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_l8_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     l8_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     l8_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := l8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- deo_param1_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_deo_param0_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_deo_param1_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_l8_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_t8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- t8_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_t8_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     t8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     t8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l533_c2_51df_return_output := t8_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- deo_param1_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_return_output := deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- l8_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_l8_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     l8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     l8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l543_c7_d631_return_output := l8_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- n8_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_n8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     n8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     n8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := n8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- deo_param0_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_deo_param0_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_deo_param1_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_l8_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_n8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l533_c2_51df_return_output;
     -- n8_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_n8_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     n8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     n8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l533_c2_51df_return_output := n8_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- deo_param0_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_return_output := deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- deo_param1_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- l8_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_l8_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     l8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     l8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := l8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- Submodule level 5
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_deo_param0_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_deo_param1_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_l8_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l533_c2_51df_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l556_c1_7044] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_return_output;

     -- deo_param1_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_return_output := deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- deo_param0_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- l8_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_l8_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     l8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     l8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l533_c2_51df_return_output := l8_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- Submodule level 6
     VAR_device_out_uxn_opcodes_h_l560_c23_82e8_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l556_c1_7044_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_deo_param0_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     REG_VAR_deo_param1 := VAR_deo_param1_MUX_uxn_opcodes_h_l533_c2_51df_return_output;
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l533_c2_51df_return_output;
     -- deo_param0_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_return_output := deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- device_out[uxn_opcodes_h_l560_c23_82e8] LATENCY=0
     -- Clock enable
     device_out_uxn_opcodes_h_l560_c23_82e8_CLOCK_ENABLE <= VAR_device_out_uxn_opcodes_h_l560_c23_82e8_CLOCK_ENABLE;
     -- Inputs
     device_out_uxn_opcodes_h_l560_c23_82e8_device_address <= VAR_device_out_uxn_opcodes_h_l560_c23_82e8_device_address;
     device_out_uxn_opcodes_h_l560_c23_82e8_value <= VAR_device_out_uxn_opcodes_h_l560_c23_82e8_value;
     device_out_uxn_opcodes_h_l560_c23_82e8_phase <= VAR_device_out_uxn_opcodes_h_l560_c23_82e8_phase;
     device_out_uxn_opcodes_h_l560_c23_82e8_previous_device_ram_read <= VAR_device_out_uxn_opcodes_h_l560_c23_82e8_previous_device_ram_read;
     device_out_uxn_opcodes_h_l560_c23_82e8_previous_ram_read <= VAR_device_out_uxn_opcodes_h_l560_c23_82e8_previous_ram_read;
     -- Outputs
     VAR_device_out_uxn_opcodes_h_l560_c23_82e8_return_output := device_out_uxn_opcodes_h_l560_c23_82e8_return_output;

     -- Submodule level 7
     REG_VAR_deo_param0 := VAR_deo_param0_MUX_uxn_opcodes_h_l533_c2_51df_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_device_out_uxn_opcodes_h_l560_c23_82e8_return_output;
     -- CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d[uxn_opcodes_h_l561_c32_e0b2] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l561_c32_e0b2_return_output := VAR_device_out_uxn_opcodes_h_l560_c23_82e8_return_output.is_device_ram_write;

     -- CONST_REF_RD_uint32_t_device_out_result_t_vram_address_d41d[uxn_opcodes_h_l565_c25_61d4] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_device_out_result_t_vram_address_d41d_uxn_opcodes_h_l565_c25_61d4_return_output := VAR_device_out_uxn_opcodes_h_l560_c23_82e8_return_output.vram_address;

     -- CONST_REF_RD_uint16_t_device_out_result_t_ram_address_d41d[uxn_opcodes_h_l566_c22_dca3] LATENCY=0
     VAR_CONST_REF_RD_uint16_t_device_out_result_t_ram_address_d41d_uxn_opcodes_h_l566_c22_dca3_return_output := VAR_device_out_uxn_opcodes_h_l560_c23_82e8_return_output.ram_address;

     -- CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d[uxn_opcodes_h_l562_c31_8d15] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l562_c31_8d15_return_output := VAR_device_out_uxn_opcodes_h_l560_c23_82e8_return_output.device_ram_address;

     -- device_out_result_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_return_output := device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d[uxn_opcodes_h_l564_c29_faf0] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l564_c29_faf0_return_output := VAR_device_out_uxn_opcodes_h_l560_c23_82e8_return_output.vram_write_layer;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d[uxn_opcodes_h_l563_c26_a98f] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l563_c26_a98f_return_output := VAR_device_out_uxn_opcodes_h_l560_c23_82e8_return_output.is_vram_write;

     -- CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d[uxn_opcodes_h_l567_c21_c2b2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l567_c21_c2b2_return_output := VAR_device_out_uxn_opcodes_h_l560_c23_82e8_return_output.u8_value;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l568_l569_DUPLICATE_6038 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l568_l569_DUPLICATE_6038_return_output := VAR_device_out_uxn_opcodes_h_l560_c23_82e8_return_output.is_deo_done;

     -- Submodule level 8
     VAR_result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_CONST_REF_RD_uint16_t_device_out_result_t_ram_address_d41d_uxn_opcodes_h_l566_c22_dca3_return_output;
     VAR_BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_left := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l568_l569_DUPLICATE_6038_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_cond := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l568_l569_DUPLICATE_6038_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_cond := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l568_l569_DUPLICATE_6038_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l561_c32_e0b2_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l563_c26_a98f_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l564_c29_faf0_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_CONST_REF_RD_uint32_t_device_out_result_t_vram_address_d41d_uxn_opcodes_h_l565_c25_61d4_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l562_c31_8d15_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l567_c21_c2b2_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_device_out_result_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     -- result_vram_address_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output := result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- device_out_result_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output := result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output := result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l568_c24_9a70] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_left;
     BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_return_output := BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_return_output;

     -- is_second_deo_MUX[uxn_opcodes_h_l569_c3_57f7] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_cond;
     is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_return_output := is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- current_deo_phase_MUX[uxn_opcodes_h_l569_c3_57f7] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_return_output := current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- Submodule level 9
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_BIN_OP_AND_uxn_opcodes_h_l568_c24_9a70_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_current_deo_phase_MUX_uxn_opcodes_h_l569_c3_57f7_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_device_out_result_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_iffalse := VAR_is_second_deo_MUX_uxn_opcodes_h_l569_c3_57f7_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_result_is_vram_write_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_result_vram_address_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- result_vram_address_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- current_deo_phase_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_return_output := current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- device_out_result_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_return_output := device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- is_second_deo_MUX[uxn_opcodes_h_l550_c7_c749] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_cond;
     is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_return_output := is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- Submodule level 10
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_current_deo_phase_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_device_out_result_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_is_second_deo_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l550_c7_c749_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_result_is_vram_write_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_result_vram_address_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- current_deo_phase_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output := result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- is_second_deo_MUX[uxn_opcodes_h_l547_c7_f1ac] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_cond;
     is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output := is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;

     -- device_out_result_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- result_vram_address_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output := result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output := result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- Submodule level 11
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_current_deo_phase_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_device_out_result_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_is_second_deo_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l547_c7_f1ac_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_result_is_vram_write_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_result_vram_address_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- result_vram_address_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- device_out_result_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_return_output := device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- is_second_deo_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_return_output := is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- current_deo_phase_MUX[uxn_opcodes_h_l543_c7_d631] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_return_output := current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_return_output;

     -- Submodule level 12
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_current_deo_phase_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     REG_VAR_device_out_result := VAR_device_out_result_MUX_uxn_opcodes_h_l533_c2_51df_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_is_second_deo_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l543_c7_d631_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_result_is_vram_write_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_result_vram_address_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output := result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output := result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- is_second_deo_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- result_vram_address_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output := result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- current_deo_phase_MUX[uxn_opcodes_h_l540_c7_7e3c] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output := current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;

     -- Submodule level 13
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_current_deo_phase_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_is_second_deo_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l540_c7_7e3c_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- is_second_deo_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_return_output := is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- current_deo_phase_MUX[uxn_opcodes_h_l533_c2_51df] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_return_output := current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_return_output;

     -- Submodule level 14
     REG_VAR_current_deo_phase := VAR_current_deo_phase_MUX_uxn_opcodes_h_l533_c2_51df_return_output;
     REG_VAR_is_second_deo := VAR_is_second_deo_MUX_uxn_opcodes_h_l533_c2_51df_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e309_uxn_opcodes_h_l577_l527_DUPLICATE_9675 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e309_uxn_opcodes_h_l577_l527_DUPLICATE_9675_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e309(
     result,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
     VAR_result_vram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l533_c2_51df_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l533_c2_51df_return_output);

     -- Submodule level 15
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e309_uxn_opcodes_h_l577_l527_DUPLICATE_9675_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e309_uxn_opcodes_h_l577_l527_DUPLICATE_9675_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_current_deo_phase <= REG_VAR_current_deo_phase;
REG_COMB_deo_param0 <= REG_VAR_deo_param0;
REG_COMB_deo_param1 <= REG_VAR_deo_param1;
REG_COMB_is_second_deo <= REG_VAR_is_second_deo;
REG_COMB_result <= REG_VAR_result;
REG_COMB_device_out_result <= REG_VAR_device_out_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     current_deo_phase <= REG_COMB_current_deo_phase;
     deo_param0 <= REG_COMB_deo_param0;
     deo_param1 <= REG_COMB_deo_param1;
     is_second_deo <= REG_COMB_is_second_deo;
     result <= REG_COMB_result;
     device_out_result <= REG_COMB_device_out_result;
 end if;
 end if;
end process;

end arch;
