-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity and_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end and_0CLK_bacf6a1d;
architecture arch of and_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l877_c6_09cd]
signal BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l877_c1_e0c4]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l877_c2_794b]
signal t8_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l877_c2_794b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l877_c2_794b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l877_c2_794b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l877_c2_794b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l877_c2_794b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l877_c2_794b]
signal result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l877_c2_794b]
signal n8_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l878_c3_efcf[uxn_opcodes_h_l878_c3_efcf]
signal printf_uxn_opcodes_h_l878_c3_efcf_uxn_opcodes_h_l878_c3_efcf_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l882_c11_f813]
signal BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l882_c7_e0ef]
signal t8_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l882_c7_e0ef]
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l882_c7_e0ef]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l882_c7_e0ef]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l882_c7_e0ef]
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l882_c7_e0ef]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l882_c7_e0ef]
signal result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l882_c7_e0ef]
signal n8_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l885_c11_d0e7]
signal BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l885_c7_e398]
signal t8_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l885_c7_e398]
signal result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l885_c7_e398]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l885_c7_e398]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l885_c7_e398]
signal result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l885_c7_e398]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l885_c7_e398]
signal result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l885_c7_e398]
signal n8_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l888_c11_ac15]
signal BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l888_c7_b980]
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l888_c7_b980]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l888_c7_b980]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l888_c7_b980]
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l888_c7_b980]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l888_c7_b980]
signal result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l888_c7_b980]
signal n8_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l888_c7_b980_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l891_c30_0a4b]
signal sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_return_output : signed(3 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l894_c21_6aee]
signal BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l896_c11_8093]
signal BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l896_c7_6126]
signal result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l896_c7_6126]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l896_c7_6126]
signal result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8c29( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd
BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_left,
BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_right,
BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_return_output);

-- t8_MUX_uxn_opcodes_h_l877_c2_794b
t8_MUX_uxn_opcodes_h_l877_c2_794b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l877_c2_794b_cond,
t8_MUX_uxn_opcodes_h_l877_c2_794b_iftrue,
t8_MUX_uxn_opcodes_h_l877_c2_794b_iffalse,
t8_MUX_uxn_opcodes_h_l877_c2_794b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b
result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_cond,
result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_return_output);

-- n8_MUX_uxn_opcodes_h_l877_c2_794b
n8_MUX_uxn_opcodes_h_l877_c2_794b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l877_c2_794b_cond,
n8_MUX_uxn_opcodes_h_l877_c2_794b_iftrue,
n8_MUX_uxn_opcodes_h_l877_c2_794b_iffalse,
n8_MUX_uxn_opcodes_h_l877_c2_794b_return_output);

-- printf_uxn_opcodes_h_l878_c3_efcf_uxn_opcodes_h_l878_c3_efcf
printf_uxn_opcodes_h_l878_c3_efcf_uxn_opcodes_h_l878_c3_efcf : entity work.printf_uxn_opcodes_h_l878_c3_efcf_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l878_c3_efcf_uxn_opcodes_h_l878_c3_efcf_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813
BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_left,
BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_right,
BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output);

-- t8_MUX_uxn_opcodes_h_l882_c7_e0ef
t8_MUX_uxn_opcodes_h_l882_c7_e0ef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l882_c7_e0ef_cond,
t8_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue,
t8_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse,
t8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef
result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_cond,
result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output);

-- n8_MUX_uxn_opcodes_h_l882_c7_e0ef
n8_MUX_uxn_opcodes_h_l882_c7_e0ef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l882_c7_e0ef_cond,
n8_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue,
n8_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse,
n8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7
BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_left,
BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_right,
BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output);

-- t8_MUX_uxn_opcodes_h_l885_c7_e398
t8_MUX_uxn_opcodes_h_l885_c7_e398 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l885_c7_e398_cond,
t8_MUX_uxn_opcodes_h_l885_c7_e398_iftrue,
t8_MUX_uxn_opcodes_h_l885_c7_e398_iffalse,
t8_MUX_uxn_opcodes_h_l885_c7_e398_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398
result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_cond,
result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_return_output);

-- n8_MUX_uxn_opcodes_h_l885_c7_e398
n8_MUX_uxn_opcodes_h_l885_c7_e398 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l885_c7_e398_cond,
n8_MUX_uxn_opcodes_h_l885_c7_e398_iftrue,
n8_MUX_uxn_opcodes_h_l885_c7_e398_iffalse,
n8_MUX_uxn_opcodes_h_l885_c7_e398_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15
BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_left,
BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_right,
BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980
result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_cond,
result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_return_output);

-- n8_MUX_uxn_opcodes_h_l888_c7_b980
n8_MUX_uxn_opcodes_h_l888_c7_b980 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l888_c7_b980_cond,
n8_MUX_uxn_opcodes_h_l888_c7_b980_iftrue,
n8_MUX_uxn_opcodes_h_l888_c7_b980_iffalse,
n8_MUX_uxn_opcodes_h_l888_c7_b980_return_output);

-- sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b
sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_ins,
sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_x,
sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_y,
sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee
BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_left,
BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_right,
BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093
BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_left,
BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_right,
BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_return_output,
 t8_MUX_uxn_opcodes_h_l877_c2_794b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_return_output,
 n8_MUX_uxn_opcodes_h_l877_c2_794b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output,
 t8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output,
 n8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output,
 t8_MUX_uxn_opcodes_h_l885_c7_e398_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_return_output,
 n8_MUX_uxn_opcodes_h_l885_c7_e398_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_return_output,
 n8_MUX_uxn_opcodes_h_l888_c7_b980_return_output,
 sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_return_output,
 BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l879_c3_2497 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c2_794b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c2_794b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c2_794b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c2_794b_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l878_c3_efcf_uxn_opcodes_h_l878_c3_efcf_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l883_c3_982e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l885_c7_e398_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l882_c7_e0ef_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l885_c7_e398_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l885_c7_e398_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l888_c7_b980_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l885_c7_e398_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l893_c3_ecea : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l888_c7_b980_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l888_c7_b980_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l888_c7_b980_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_e70a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_ed0c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_ab19_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_7a42_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l888_l882_l896_l885_DUPLICATE_c0be_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l888_l885_DUPLICATE_8f88_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l902_l873_DUPLICATE_dc8c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l883_c3_982e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l883_c3_982e;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l879_c3_2497 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l879_c3_2497;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l893_c3_ecea := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l893_c3_ecea;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_y := resize(to_signed(-1, 2), 4);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l877_c2_794b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l885_c7_e398_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l888_c7_b980_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_left := VAR_phase;
     VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l888_c7_b980_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l885_c7_e398_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l877_c2_794b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l885_c7_e398_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l877_c6_09cd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_left;
     BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output := BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l888_c11_ac15] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_left;
     BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_return_output := BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l885_c11_d0e7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_left;
     BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output := BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l891_c30_0a4b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_ins;
     sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_x;
     sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_return_output := sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_7a42 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_7a42_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_ed0c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_ed0c_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l882_c11_f813] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_left;
     BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output := BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l894_c21_6aee] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_left;
     BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_return_output := BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_e70a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_e70a_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l888_l885_DUPLICATE_8f88 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l888_l885_DUPLICATE_8f88_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_ab19 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_ab19_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l888_l882_l896_l885_DUPLICATE_c0be LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l888_l882_l896_l885_DUPLICATE_c0be_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l896_c11_8093] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_left;
     BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_return_output := BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_return_output;

     -- Submodule level 1
     VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_iftrue := VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_6aee_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l877_c2_794b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l877_c2_794b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_09cd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l882_c7_e0ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l882_c7_e0ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_f813_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l885_c7_e398_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l885_c7_e398_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_d0e7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l888_c7_b980_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_ac15_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_8093_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_ab19_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_ab19_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_ab19_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_ab19_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l888_l882_l896_l885_DUPLICATE_c0be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l888_l882_l896_l885_DUPLICATE_c0be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l888_l882_l896_l885_DUPLICATE_c0be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l888_l882_l896_l885_DUPLICATE_c0be_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_e70a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_e70a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_e70a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_e70a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_ed0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_ed0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_ed0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l877_l882_l896_l885_DUPLICATE_ed0c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l888_l885_DUPLICATE_8f88_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l888_l885_DUPLICATE_8f88_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_7a42_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_7a42_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_7a42_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l877_l888_l882_l885_DUPLICATE_7a42_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0a4b_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l877_c1_e0c4] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l896_c7_6126] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l888_c7_b980] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l888_c7_b980] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l888_c7_b980] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_cond;
     result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_return_output := result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l896_c7_6126] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_return_output;

     -- t8_MUX[uxn_opcodes_h_l885_c7_e398] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l885_c7_e398_cond <= VAR_t8_MUX_uxn_opcodes_h_l885_c7_e398_cond;
     t8_MUX_uxn_opcodes_h_l885_c7_e398_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l885_c7_e398_iftrue;
     t8_MUX_uxn_opcodes_h_l885_c7_e398_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l885_c7_e398_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l885_c7_e398_return_output := t8_MUX_uxn_opcodes_h_l885_c7_e398_return_output;

     -- n8_MUX[uxn_opcodes_h_l888_c7_b980] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l888_c7_b980_cond <= VAR_n8_MUX_uxn_opcodes_h_l888_c7_b980_cond;
     n8_MUX_uxn_opcodes_h_l888_c7_b980_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l888_c7_b980_iftrue;
     n8_MUX_uxn_opcodes_h_l888_c7_b980_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l888_c7_b980_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l888_c7_b980_return_output := n8_MUX_uxn_opcodes_h_l888_c7_b980_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l896_c7_6126] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l878_c3_efcf_uxn_opcodes_h_l878_c3_efcf_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_e0c4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l885_c7_e398_iffalse := VAR_n8_MUX_uxn_opcodes_h_l888_c7_b980_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_6126_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_6126_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_6126_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_b980_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_b980_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse := VAR_t8_MUX_uxn_opcodes_h_l885_c7_e398_return_output;
     -- printf_uxn_opcodes_h_l878_c3_efcf[uxn_opcodes_h_l878_c3_efcf] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l878_c3_efcf_uxn_opcodes_h_l878_c3_efcf_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l878_c3_efcf_uxn_opcodes_h_l878_c3_efcf_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l885_c7_e398] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l888_c7_b980] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l888_c7_b980] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l888_c7_b980] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_return_output;

     -- t8_MUX[uxn_opcodes_h_l882_c7_e0ef] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l882_c7_e0ef_cond <= VAR_t8_MUX_uxn_opcodes_h_l882_c7_e0ef_cond;
     t8_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue;
     t8_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output := t8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;

     -- n8_MUX[uxn_opcodes_h_l885_c7_e398] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l885_c7_e398_cond <= VAR_n8_MUX_uxn_opcodes_h_l885_c7_e398_cond;
     n8_MUX_uxn_opcodes_h_l885_c7_e398_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l885_c7_e398_iftrue;
     n8_MUX_uxn_opcodes_h_l885_c7_e398_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l885_c7_e398_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l885_c7_e398_return_output := n8_MUX_uxn_opcodes_h_l885_c7_e398_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l885_c7_e398] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_cond;
     result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_return_output := result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l885_c7_e398] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse := VAR_n8_MUX_uxn_opcodes_h_l885_c7_e398_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_b980_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_b980_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_b980_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_e398_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_e398_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l877_c2_794b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l885_c7_e398] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l882_c7_e0ef] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_cond;
     result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output := result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l885_c7_e398] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_return_output;

     -- t8_MUX[uxn_opcodes_h_l877_c2_794b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l877_c2_794b_cond <= VAR_t8_MUX_uxn_opcodes_h_l877_c2_794b_cond;
     t8_MUX_uxn_opcodes_h_l877_c2_794b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l877_c2_794b_iftrue;
     t8_MUX_uxn_opcodes_h_l877_c2_794b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l877_c2_794b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l877_c2_794b_return_output := t8_MUX_uxn_opcodes_h_l877_c2_794b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l885_c7_e398] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l882_c7_e0ef] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;

     -- n8_MUX[uxn_opcodes_h_l882_c7_e0ef] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l882_c7_e0ef_cond <= VAR_n8_MUX_uxn_opcodes_h_l882_c7_e0ef_cond;
     n8_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue;
     n8_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output := n8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l882_c7_e0ef] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l877_c2_794b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_e398_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_e398_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_e398_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l877_c2_794b_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l882_c7_e0ef] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l877_c2_794b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l877_c2_794b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_return_output := result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l882_c7_e0ef] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;

     -- n8_MUX[uxn_opcodes_h_l877_c2_794b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l877_c2_794b_cond <= VAR_n8_MUX_uxn_opcodes_h_l877_c2_794b_cond;
     n8_MUX_uxn_opcodes_h_l877_c2_794b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l877_c2_794b_iftrue;
     n8_MUX_uxn_opcodes_h_l877_c2_794b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l877_c2_794b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l877_c2_794b_return_output := n8_MUX_uxn_opcodes_h_l877_c2_794b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l877_c2_794b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l882_c7_e0ef] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l877_c2_794b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_e0ef_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l877_c2_794b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l877_c2_794b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l877_c2_794b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l902_l873_DUPLICATE_dc8c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l902_l873_DUPLICATE_dc8c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8c29(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_794b_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_794b_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_794b_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_794b_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_794b_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l902_l873_DUPLICATE_dc8c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l902_l873_DUPLICATE_dc8c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
