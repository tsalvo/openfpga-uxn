-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 50
entity mul_0CLK_fedec265 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end mul_0CLK_fedec265;
architecture arch of mul_0CLK_fedec265 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2095_c6_a51c]
signal BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2095_c2_fe4c]
signal n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2095_c2_fe4c]
signal t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2095_c2_fe4c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2095_c2_fe4c]
signal result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2095_c2_fe4c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2095_c2_fe4c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2095_c2_fe4c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2095_c2_fe4c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2100_c11_26f4]
signal BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2100_c7_eef8]
signal n8_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2100_c7_eef8]
signal t8_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2100_c7_eef8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2100_c7_eef8]
signal result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2100_c7_eef8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2100_c7_eef8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2100_c7_eef8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2100_c7_eef8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2103_c11_4818]
signal BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2103_c7_1bb7]
signal n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2103_c7_1bb7]
signal t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2103_c7_1bb7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2103_c7_1bb7]
signal result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2103_c7_1bb7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2103_c7_1bb7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2103_c7_1bb7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2103_c7_1bb7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2107_c11_3139]
signal BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2107_c7_421b]
signal n8_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2107_c7_421b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2107_c7_421b]
signal result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2107_c7_421b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2107_c7_421b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2107_c7_421b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2107_c7_421b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2110_c11_34ec]
signal BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2110_c7_fce2]
signal n8_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2110_c7_fce2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2110_c7_fce2]
signal result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2110_c7_fce2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2110_c7_fce2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2110_c7_fce2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2110_c7_fce2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2113_c30_ebf1]
signal sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_return_output : signed(3 downto 0);

-- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l2116_c21_d4c5]
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_left : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_right : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2118_c11_4c6f]
signal BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2118_c7_b0ac]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2118_c7_b0ac]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2118_c7_b0ac]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_3345( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c
BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_left,
BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_right,
BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output);

-- n8_MUX_uxn_opcodes_h_l2095_c2_fe4c
n8_MUX_uxn_opcodes_h_l2095_c2_fe4c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond,
n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue,
n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse,
n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output);

-- t8_MUX_uxn_opcodes_h_l2095_c2_fe4c
t8_MUX_uxn_opcodes_h_l2095_c2_fe4c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond,
t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue,
t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse,
t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c
result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c
result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c
result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c
result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4
BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_left,
BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_right,
BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output);

-- n8_MUX_uxn_opcodes_h_l2100_c7_eef8
n8_MUX_uxn_opcodes_h_l2100_c7_eef8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2100_c7_eef8_cond,
n8_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue,
n8_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse,
n8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output);

-- t8_MUX_uxn_opcodes_h_l2100_c7_eef8
t8_MUX_uxn_opcodes_h_l2100_c7_eef8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2100_c7_eef8_cond,
t8_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue,
t8_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse,
t8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8
result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8
result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8
result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8
result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818
BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_left,
BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_right,
BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output);

-- n8_MUX_uxn_opcodes_h_l2103_c7_1bb7
n8_MUX_uxn_opcodes_h_l2103_c7_1bb7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond,
n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue,
n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse,
n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output);

-- t8_MUX_uxn_opcodes_h_l2103_c7_1bb7
t8_MUX_uxn_opcodes_h_l2103_c7_1bb7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond,
t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue,
t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse,
t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7
result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond,
result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7
result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7
result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7
result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7
result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139
BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_left,
BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_right,
BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_return_output);

-- n8_MUX_uxn_opcodes_h_l2107_c7_421b
n8_MUX_uxn_opcodes_h_l2107_c7_421b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2107_c7_421b_cond,
n8_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue,
n8_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse,
n8_MUX_uxn_opcodes_h_l2107_c7_421b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b
result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b
result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b
result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b
result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec
BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_left,
BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_right,
BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_return_output);

-- n8_MUX_uxn_opcodes_h_l2110_c7_fce2
n8_MUX_uxn_opcodes_h_l2110_c7_fce2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2110_c7_fce2_cond,
n8_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue,
n8_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse,
n8_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2
result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2
result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2
result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2
result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1
sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_ins,
sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_x,
sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_y,
sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_return_output);

-- BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5 : entity work.BIN_OP_INFERRED_MULT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_left,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_right,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f
BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_left,
BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_right,
BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac
result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac
result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac
result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output,
 n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output,
 t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output,
 n8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output,
 t8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output,
 n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output,
 t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_return_output,
 n8_MUX_uxn_opcodes_h_l2107_c7_421b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_return_output,
 n8_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output,
 sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_return_output,
 BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2097_c3_4817 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2101_c3_a8df : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2105_c3_7428 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2108_c3_0732 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2115_c3_ca3e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2110_c7_fce2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l2116_c3_aa4a : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_bb7c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_dcc5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_f246_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_b7dd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2118_l2110_l2107_l2103_l2100_DUPLICATE_b629_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2124_l2091_DUPLICATE_9cc4_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2108_c3_0732 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2108_c3_0732;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2115_c3_ca3e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2115_c3_ca3e;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_right := to_unsigned(5, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2101_c3_a8df := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2101_c3_a8df;
     VAR_sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2097_c3_4817 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2097_c3_4817;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2105_c3_7428 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2105_c3_7428;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_left := VAR_phase;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2100_c11_26f4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_dcc5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_dcc5_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2107_c11_3139] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_left;
     BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_return_output := BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2118_c11_4c6f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2118_l2110_l2107_l2103_l2100_DUPLICATE_b629 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2118_l2110_l2107_l2103_l2100_DUPLICATE_b629_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2103_c11_4818] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_left;
     BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output := BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2095_c6_a51c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output;

     -- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l2116_c21_d4c5] LATENCY=0
     -- Inputs
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_left <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_left;
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_right <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_right;
     -- Outputs
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_return_output := BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_bb7c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_bb7c_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_b7dd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_b7dd_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2110_c11_34ec] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_left;
     BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_return_output := BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2110_c7_fce2] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2110_c7_fce2_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_f246 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_f246_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l2113_c30_ebf1] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_ins;
     sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_x;
     sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_return_output := sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2095_c6_a51c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2100_c7_eef8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2100_c7_eef8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_26f4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2103_c11_4818_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2107_c7_421b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_3139_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2110_c7_fce2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2110_c11_34ec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2118_c11_4c6f_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l2116_c3_aa4a := resize(VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2116_c21_d4c5_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_f246_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_f246_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_f246_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_f246_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_f246_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2118_l2110_l2107_l2103_l2100_DUPLICATE_b629_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2118_l2110_l2107_l2103_l2100_DUPLICATE_b629_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2118_l2110_l2107_l2103_l2100_DUPLICATE_b629_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2118_l2110_l2107_l2103_l2100_DUPLICATE_b629_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2118_l2110_l2107_l2103_l2100_DUPLICATE_b629_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_b7dd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_b7dd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_b7dd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_b7dd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_b7dd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_dcc5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_dcc5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_dcc5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_dcc5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2118_l2107_l2103_l2100_l2095_DUPLICATE_dcc5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_bb7c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_bb7c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_bb7c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_bb7c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2110_l2107_l2103_l2100_l2095_DUPLICATE_bb7c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2110_c7_fce2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2113_c30_ebf1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue := VAR_result_u8_value_uxn_opcodes_h_l2116_c3_aa4a;
     -- t8_MUX[uxn_opcodes_h_l2103_c7_1bb7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond <= VAR_t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond;
     t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue;
     t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output := t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;

     -- n8_MUX[uxn_opcodes_h_l2110_c7_fce2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2110_c7_fce2_cond <= VAR_n8_MUX_uxn_opcodes_h_l2110_c7_fce2_cond;
     n8_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue;
     n8_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output := n8_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2110_c7_fce2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2118_c7_b0ac] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2118_c7_b0ac] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2118_c7_b0ac] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2110_c7_fce2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2110_c7_fce2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2118_c7_b0ac_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2107_c7_421b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2107_c7_421b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2110_c7_fce2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;

     -- n8_MUX[uxn_opcodes_h_l2107_c7_421b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2107_c7_421b_cond <= VAR_n8_MUX_uxn_opcodes_h_l2107_c7_421b_cond;
     n8_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue;
     n8_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2107_c7_421b_return_output := n8_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;

     -- t8_MUX[uxn_opcodes_h_l2100_c7_eef8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2100_c7_eef8_cond <= VAR_t8_MUX_uxn_opcodes_h_l2100_c7_eef8_cond;
     t8_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue;
     t8_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output := t8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2107_c7_421b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2110_c7_fce2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2110_c7_fce2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2110_c7_fce2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2103_c7_1bb7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;

     -- t8_MUX[uxn_opcodes_h_l2095_c2_fe4c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond <= VAR_t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond;
     t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue;
     t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output := t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2103_c7_1bb7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output := result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2107_c7_421b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2103_c7_1bb7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;

     -- n8_MUX[uxn_opcodes_h_l2103_c7_1bb7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond <= VAR_n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond;
     n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue;
     n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output := n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2107_c7_421b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2107_c7_421b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_421b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2103_c7_1bb7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2100_c7_eef8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2100_c7_eef8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2103_c7_1bb7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2103_c7_1bb7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;

     -- n8_MUX[uxn_opcodes_h_l2100_c7_eef8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2100_c7_eef8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2100_c7_eef8_cond;
     n8_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue;
     n8_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output := n8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2100_c7_eef8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2103_c7_1bb7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2100_c7_eef8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;

     -- n8_MUX[uxn_opcodes_h_l2095_c2_fe4c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond;
     n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue;
     n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output := n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2095_c2_fe4c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2095_c2_fe4c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2100_c7_eef8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2095_c2_fe4c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2100_c7_eef8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_eef8_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2095_c2_fe4c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2095_c2_fe4c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2095_c2_fe4c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2124_l2091_DUPLICATE_9cc4 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2124_l2091_DUPLICATE_9cc4_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3345(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2095_c2_fe4c_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2124_l2091_DUPLICATE_9cc4_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2124_l2091_DUPLICATE_9cc4_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
