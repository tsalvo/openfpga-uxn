-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity neq_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_226c8821;
architecture arch of neq_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1265_c6_30ef]
signal BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1265_c2_8488]
signal t8_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1265_c2_8488]
signal n8_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1265_c2_8488]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1265_c2_8488]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1265_c2_8488]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1265_c2_8488]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1265_c2_8488]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1265_c2_8488]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1265_c2_8488]
signal result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1265_c2_8488]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1265_c2_8488]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1278_c11_34d5]
signal BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1278_c7_0ddd]
signal t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1278_c7_0ddd]
signal n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1278_c7_0ddd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1278_c7_0ddd]
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1278_c7_0ddd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1278_c7_0ddd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1278_c7_0ddd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1281_c11_0e6a]
signal BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1281_c7_7f25]
signal t8_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1281_c7_7f25]
signal n8_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1281_c7_7f25]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1281_c7_7f25]
signal result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1281_c7_7f25]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1281_c7_7f25]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1281_c7_7f25]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1284_c11_8e20]
signal BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1284_c7_6005]
signal n8_MUX_uxn_opcodes_h_l1284_c7_6005_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1284_c7_6005_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1284_c7_6005]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1284_c7_6005]
signal result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1284_c7_6005]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1284_c7_6005]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1284_c7_6005]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1286_c30_1029]
signal sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1289_c21_171b]
signal BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1289_c21_df63]
signal MUX_uxn_opcodes_h_l1289_c21_df63_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1289_c21_df63_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1289_c21_df63_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1289_c21_df63_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef
BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_left,
BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_right,
BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output);

-- t8_MUX_uxn_opcodes_h_l1265_c2_8488
t8_MUX_uxn_opcodes_h_l1265_c2_8488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1265_c2_8488_cond,
t8_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue,
t8_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse,
t8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output);

-- n8_MUX_uxn_opcodes_h_l1265_c2_8488
n8_MUX_uxn_opcodes_h_l1265_c2_8488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1265_c2_8488_cond,
n8_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue,
n8_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse,
n8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488
result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488
result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488
result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488
result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488
result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488
result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_cond,
result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488
result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_left,
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_right,
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_return_output);

-- t8_MUX_uxn_opcodes_h_l1278_c7_0ddd
t8_MUX_uxn_opcodes_h_l1278_c7_0ddd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond,
t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue,
t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse,
t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output);

-- n8_MUX_uxn_opcodes_h_l1278_c7_0ddd
n8_MUX_uxn_opcodes_h_l1278_c7_0ddd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond,
n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue,
n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse,
n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond,
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a
BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_left,
BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_right,
BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_return_output);

-- t8_MUX_uxn_opcodes_h_l1281_c7_7f25
t8_MUX_uxn_opcodes_h_l1281_c7_7f25 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1281_c7_7f25_cond,
t8_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue,
t8_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse,
t8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output);

-- n8_MUX_uxn_opcodes_h_l1281_c7_7f25
n8_MUX_uxn_opcodes_h_l1281_c7_7f25 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1281_c7_7f25_cond,
n8_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue,
n8_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse,
n8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25
result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25
result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_cond,
result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25
result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25
result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20
BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_left,
BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_right,
BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_return_output);

-- n8_MUX_uxn_opcodes_h_l1284_c7_6005
n8_MUX_uxn_opcodes_h_l1284_c7_6005 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1284_c7_6005_cond,
n8_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue,
n8_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse,
n8_MUX_uxn_opcodes_h_l1284_c7_6005_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005
result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_cond,
result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005
result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1286_c30_1029
sp_relative_shift_uxn_opcodes_h_l1286_c30_1029 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_ins,
sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_x,
sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_y,
sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b
BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_left,
BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_right,
BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_return_output);

-- MUX_uxn_opcodes_h_l1289_c21_df63
MUX_uxn_opcodes_h_l1289_c21_df63 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1289_c21_df63_cond,
MUX_uxn_opcodes_h_l1289_c21_df63_iftrue,
MUX_uxn_opcodes_h_l1289_c21_df63_iffalse,
MUX_uxn_opcodes_h_l1289_c21_df63_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output,
 t8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
 n8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_return_output,
 t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output,
 n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_return_output,
 t8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output,
 n8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_return_output,
 n8_MUX_uxn_opcodes_h_l1284_c7_6005_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_return_output,
 sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_return_output,
 MUX_uxn_opcodes_h_l1289_c21_df63_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1270_c3_d394 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1275_c3_4825 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1279_c3_0e72 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1284_c7_6005_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1284_c7_6005_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1288_c3_3266 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1289_c21_df63_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1289_c21_df63_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1289_c21_df63_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1289_c21_df63_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1265_l1284_l1278_l1281_DUPLICATE_4b04_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_fde9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_d6b9_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_fcb9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1284_l1281_DUPLICATE_c792_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1293_l1261_DUPLICATE_1189_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1289_c21_df63_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1288_c3_3266 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1288_c3_3266;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1279_c3_0e72 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1279_c3_0e72;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1270_c3_d394 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1270_c3_d394;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1275_c3_4825 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1275_c3_4825;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_right := to_unsigned(2, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1289_c21_df63_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse := t8;
     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1265_c2_8488_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1289_c21_171b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1265_c2_8488_return_output := result.is_stack_index_flipped;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1265_c2_8488_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1278_c11_34d5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1284_c11_8e20] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_left;
     BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_return_output := BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1286_c30_1029] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_ins;
     sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_x;
     sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_return_output := sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_fde9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_fde9_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1265_l1284_l1278_l1281_DUPLICATE_4b04 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1265_l1284_l1278_l1281_DUPLICATE_4b04_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_fcb9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_fcb9_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1284_l1281_DUPLICATE_c792 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1284_l1281_DUPLICATE_c792_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1281_c11_0e6a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1265_c6_30ef] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_left;
     BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output := BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_d6b9 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_d6b9_return_output := result.sp_relative_shift;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1265_c2_8488_return_output := result.is_vram_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1265_c2_8488_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1265_c2_8488_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1265_c6_30ef_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_34d5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1281_c7_7f25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1281_c7_7f25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1281_c11_0e6a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1284_c7_6005_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_8e20_return_output;
     VAR_MUX_uxn_opcodes_h_l1289_c21_df63_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1289_c21_171b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_d6b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_d6b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_d6b9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_fde9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_fde9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_fde9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_fcb9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_fcb9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1284_l1278_l1281_DUPLICATE_fcb9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1284_l1281_DUPLICATE_c792_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1284_l1281_DUPLICATE_c792_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1265_l1284_l1278_l1281_DUPLICATE_4b04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1265_l1284_l1278_l1281_DUPLICATE_4b04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1265_l1284_l1278_l1281_DUPLICATE_4b04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1265_l1284_l1278_l1281_DUPLICATE_4b04_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1265_c2_8488_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1265_c2_8488_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1265_c2_8488_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1265_c2_8488_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1286_c30_1029_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1284_c7_6005] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1284_c7_6005] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1284_c7_6005] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1284_c7_6005] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_return_output;

     -- MUX[uxn_opcodes_h_l1289_c21_df63] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1289_c21_df63_cond <= VAR_MUX_uxn_opcodes_h_l1289_c21_df63_cond;
     MUX_uxn_opcodes_h_l1289_c21_df63_iftrue <= VAR_MUX_uxn_opcodes_h_l1289_c21_df63_iftrue;
     MUX_uxn_opcodes_h_l1289_c21_df63_iffalse <= VAR_MUX_uxn_opcodes_h_l1289_c21_df63_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1289_c21_df63_return_output := MUX_uxn_opcodes_h_l1289_c21_df63_return_output;

     -- t8_MUX[uxn_opcodes_h_l1281_c7_7f25] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1281_c7_7f25_cond <= VAR_t8_MUX_uxn_opcodes_h_l1281_c7_7f25_cond;
     t8_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue;
     t8_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output := t8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;

     -- n8_MUX[uxn_opcodes_h_l1284_c7_6005] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1284_c7_6005_cond <= VAR_n8_MUX_uxn_opcodes_h_l1284_c7_6005_cond;
     n8_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue;
     n8_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1284_c7_6005_return_output := n8_MUX_uxn_opcodes_h_l1284_c7_6005_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue := VAR_MUX_uxn_opcodes_h_l1289_c21_df63_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1284_c7_6005_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_6005_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_6005_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c7_6005_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c7_6005_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1281_c7_7f25] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1281_c7_7f25] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1284_c7_6005] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_return_output := result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_return_output;

     -- n8_MUX[uxn_opcodes_h_l1281_c7_7f25] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1281_c7_7f25_cond <= VAR_n8_MUX_uxn_opcodes_h_l1281_c7_7f25_cond;
     n8_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue;
     n8_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output := n8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1281_c7_7f25] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1281_c7_7f25] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;

     -- t8_MUX[uxn_opcodes_h_l1278_c7_0ddd] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond <= VAR_t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond;
     t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue;
     t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output := t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1284_c7_6005_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1278_c7_0ddd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1278_c7_0ddd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1278_c7_0ddd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1281_c7_7f25] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output := result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;

     -- t8_MUX[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1265_c2_8488_cond <= VAR_t8_MUX_uxn_opcodes_h_l1265_c2_8488_cond;
     t8_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue;
     t8_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output := t8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output;

     -- n8_MUX[uxn_opcodes_h_l1278_c7_0ddd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond <= VAR_n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond;
     n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue;
     n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output := n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1278_c7_0ddd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1281_c7_7f25_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_return_output;

     -- n8_MUX[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1265_c2_8488_cond <= VAR_n8_MUX_uxn_opcodes_h_l1265_c2_8488_cond;
     n8_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue;
     n8_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output := n8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1278_c7_0ddd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output := result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1265_c2_8488_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_0ddd_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1265_c2_8488] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_return_output := result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1293_l1261_DUPLICATE_1189 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1293_l1261_DUPLICATE_1189_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1265_c2_8488_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1265_c2_8488_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1293_l1261_DUPLICATE_1189_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1293_l1261_DUPLICATE_1189_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
