-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity sub1_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub1_0CLK_64d180f1;
architecture arch of sub1_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2462_c6_f81d]
signal BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2462_c2_732f]
signal n8_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2462_c2_732f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2462_c2_732f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2462_c2_732f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2462_c2_732f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2462_c2_732f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2462_c2_732f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2462_c2_732f]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2462_c2_732f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2462_c2_732f]
signal result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2462_c2_732f]
signal t8_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2475_c11_83ca]
signal BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2475_c7_3947]
signal n8_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2475_c7_3947]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2475_c7_3947]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2475_c7_3947]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2475_c7_3947]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2475_c7_3947]
signal result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2475_c7_3947]
signal t8_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2478_c11_ee64]
signal BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2478_c7_0bf1]
signal n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2478_c7_0bf1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2478_c7_0bf1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2478_c7_0bf1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2478_c7_0bf1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2478_c7_0bf1]
signal result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2478_c7_0bf1]
signal t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2481_c11_72bf]
signal BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2481_c7_481e]
signal n8_MUX_uxn_opcodes_h_l2481_c7_481e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2481_c7_481e_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2481_c7_481e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2481_c7_481e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2481_c7_481e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2481_c7_481e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2481_c7_481e]
signal result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2483_c30_695b]
signal sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_return_output : signed(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2486_c21_1118]
signal BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_04b4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d
BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_left,
BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_right,
BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output);

-- n8_MUX_uxn_opcodes_h_l2462_c2_732f
n8_MUX_uxn_opcodes_h_l2462_c2_732f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2462_c2_732f_cond,
n8_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue,
n8_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse,
n8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f
result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f
result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f
result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f
result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f
result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f
result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_return_output);

-- t8_MUX_uxn_opcodes_h_l2462_c2_732f
t8_MUX_uxn_opcodes_h_l2462_c2_732f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2462_c2_732f_cond,
t8_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue,
t8_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse,
t8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca
BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_left,
BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_right,
BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_return_output);

-- n8_MUX_uxn_opcodes_h_l2475_c7_3947
n8_MUX_uxn_opcodes_h_l2475_c7_3947 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2475_c7_3947_cond,
n8_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue,
n8_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse,
n8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947
result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947
result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947
result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947
result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_cond,
result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_return_output);

-- t8_MUX_uxn_opcodes_h_l2475_c7_3947
t8_MUX_uxn_opcodes_h_l2475_c7_3947 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2475_c7_3947_cond,
t8_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue,
t8_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse,
t8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64
BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_left,
BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_right,
BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_return_output);

-- n8_MUX_uxn_opcodes_h_l2478_c7_0bf1
n8_MUX_uxn_opcodes_h_l2478_c7_0bf1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond,
n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue,
n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse,
n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1
result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1
result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1
result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1
result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond,
result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output);

-- t8_MUX_uxn_opcodes_h_l2478_c7_0bf1
t8_MUX_uxn_opcodes_h_l2478_c7_0bf1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond,
t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue,
t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse,
t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf
BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_left,
BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_right,
BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_return_output);

-- n8_MUX_uxn_opcodes_h_l2481_c7_481e
n8_MUX_uxn_opcodes_h_l2481_c7_481e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2481_c7_481e_cond,
n8_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue,
n8_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse,
n8_MUX_uxn_opcodes_h_l2481_c7_481e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e
result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e
result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e
result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2483_c30_695b
sp_relative_shift_uxn_opcodes_h_l2483_c30_695b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_ins,
sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_x,
sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_y,
sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118
BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_left,
BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_right,
BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output,
 n8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
 t8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_return_output,
 n8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_return_output,
 t8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_return_output,
 n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output,
 t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_return_output,
 n8_MUX_uxn_opcodes_h_l2481_c7_481e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_return_output,
 sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2472_c3_1337 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2467_c3_9de3 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2462_c2_732f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2476_c3_c79b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2475_c7_3947_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2481_c7_481e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2481_c7_481e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2485_c3_f4ed : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2475_l2478_l2462_l2481_DUPLICATE_09da_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_1372_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_dc81_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_0561_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2478_l2481_DUPLICATE_40ab_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2490_l2458_DUPLICATE_a8fe_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2472_c3_1337 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2472_c3_1337;
     VAR_sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2467_c3_9de3 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2467_c3_9de3;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_right := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_right := to_unsigned(3, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2476_c3_c79b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2476_c3_c79b;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2485_c3_f4ed := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2485_c3_f4ed;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse := t8;
     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2462_c2_732f_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2462_c6_f81d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_0561 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_0561_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2478_l2481_DUPLICATE_40ab LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2478_l2481_DUPLICATE_40ab_return_output := result.stack_address_sp_offset;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2462_c2_732f_return_output := result.is_ram_write;

     -- sp_relative_shift[uxn_opcodes_h_l2483_c30_695b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_ins;
     sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_x;
     sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_return_output := sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2481_c11_72bf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_left;
     BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_return_output := BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_1372 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_1372_return_output := result.sp_relative_shift;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2462_c2_732f_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2475_l2478_l2462_l2481_DUPLICATE_09da LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2475_l2478_l2462_l2481_DUPLICATE_09da_return_output := result.u8_value;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2486_c21_1118] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2462_c2_732f_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_dc81 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_dc81_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2478_c11_ee64] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_left;
     BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_return_output := BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2475_c11_83ca] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_left;
     BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_return_output := BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2462_c2_732f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2462_c2_732f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c6_f81d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2475_c7_3947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2475_c7_3947_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2475_c11_83ca_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c11_ee64_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2481_c7_481e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2481_c11_72bf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2486_c21_1118_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_1372_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_1372_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_1372_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_dc81_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_dc81_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_dc81_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_0561_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_0561_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2475_l2478_l2481_DUPLICATE_0561_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2478_l2481_DUPLICATE_40ab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2478_l2481_DUPLICATE_40ab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2475_l2478_l2462_l2481_DUPLICATE_09da_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2475_l2478_l2462_l2481_DUPLICATE_09da_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2475_l2478_l2462_l2481_DUPLICATE_09da_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2475_l2478_l2462_l2481_DUPLICATE_09da_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2462_c2_732f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2462_c2_732f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2462_c2_732f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2462_c2_732f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2483_c30_695b_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2481_c7_481e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2481_c7_481e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2481_c7_481e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2481_c7_481e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_return_output;

     -- t8_MUX[uxn_opcodes_h_l2478_c7_0bf1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond <= VAR_t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond;
     t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue;
     t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output := t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2481_c7_481e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2481_c7_481e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2481_c7_481e_cond <= VAR_n8_MUX_uxn_opcodes_h_l2481_c7_481e_cond;
     n8_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2481_c7_481e_iftrue;
     n8_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2481_c7_481e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2481_c7_481e_return_output := n8_MUX_uxn_opcodes_h_l2481_c7_481e_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2481_c7_481e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2481_c7_481e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2481_c7_481e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2481_c7_481e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2481_c7_481e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2481_c7_481e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2478_c7_0bf1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;

     -- n8_MUX[uxn_opcodes_h_l2478_c7_0bf1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond <= VAR_n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond;
     n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue;
     n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output := n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2478_c7_0bf1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2478_c7_0bf1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2478_c7_0bf1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output := result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;

     -- t8_MUX[uxn_opcodes_h_l2475_c7_3947] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2475_c7_3947_cond <= VAR_t8_MUX_uxn_opcodes_h_l2475_c7_3947_cond;
     t8_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue;
     t8_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output := t8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2478_c7_0bf1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c7_0bf1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2475_c7_3947] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_return_output := result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2475_c7_3947] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2475_c7_3947] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;

     -- t8_MUX[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2462_c2_732f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2462_c2_732f_cond;
     t8_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue;
     t8_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output := t8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2475_c7_3947] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2475_c7_3947] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;

     -- n8_MUX[uxn_opcodes_h_l2475_c7_3947] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2475_c7_3947_cond <= VAR_n8_MUX_uxn_opcodes_h_l2475_c7_3947_cond;
     n8_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2475_c7_3947_iftrue;
     n8_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2475_c7_3947_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output := n8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2475_c7_3947_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_return_output;

     -- n8_MUX[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2462_c2_732f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2462_c2_732f_cond;
     n8_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue;
     n8_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output := n8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2462_c2_732f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2462_c2_732f_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2490_l2458_DUPLICATE_a8fe LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2490_l2458_DUPLICATE_a8fe_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_04b4(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2462_c2_732f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c2_732f_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2490_l2458_DUPLICATE_a8fe_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2490_l2458_DUPLICATE_a8fe_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
