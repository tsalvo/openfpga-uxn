-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 17
entity VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_0CLK_83e31706 is
port(
 elem_val : in unsigned(7 downto 0);
 ref_toks_0 : in uint8_t_8;
 var_dim_0 : in unsigned(2 downto 0);
 return_output : out uint8_t_array_8_t);
end VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_0CLK_83e31706;
architecture arch of VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_0CLK_83e31706 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_return_output : unsigned(0 downto 0);

-- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43]
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_cond : unsigned(0 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_iftrue : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_iffalse : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_return_output : unsigned(0 downto 0);

-- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea]
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_cond : unsigned(0 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_iftrue : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_iffalse : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_return_output : unsigned(0 downto 0);

-- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913]
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_cond : unsigned(0 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_iftrue : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_iffalse : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_return_output : unsigned(0 downto 0);

-- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412]
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_cond : unsigned(0 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_iftrue : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_iffalse : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_return_output : unsigned(0 downto 0);

-- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859]
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_cond : unsigned(0 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_iftrue : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_iffalse : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_return_output : unsigned(0 downto 0);

-- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a]
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_cond : unsigned(0 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_iftrue : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_iffalse : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_return_output : unsigned(0 downto 0);

-- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678]
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_cond : unsigned(0 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_iftrue : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_iffalse : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_return_output : unsigned(0 downto 0);

-- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531]
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_cond : unsigned(0 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_iftrue : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_iffalse : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_return_output : unsigned(7 downto 0);

function CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_e759( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return uint8_t_array_8_t is
 
  variable base : uint8_t_array_8_t; 
  variable return_output : uint8_t_array_8_t;
begin
      base.data(2) := ref_toks_0;
      base.data(5) := ref_toks_1;
      base.data(1) := ref_toks_2;
      base.data(4) := ref_toks_3;
      base.data(7) := ref_toks_4;
      base.data(0) := ref_toks_5;
      base.data(6) := ref_toks_6;
      base.data(3) := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8 : entity work.BIN_OP_EQ_uint3_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_return_output);

-- rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_cond,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_iftrue,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_iffalse,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_return_output);

-- rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_cond,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_iftrue,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_iffalse,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15 : entity work.BIN_OP_EQ_uint3_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_return_output);

-- rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_cond,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_iftrue,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_iffalse,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_return_output);

-- rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_cond,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_iftrue,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_iffalse,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7 : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_return_output);

-- rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_cond,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_iftrue,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_iffalse,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46 : entity work.BIN_OP_EQ_uint3_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_return_output);

-- rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_cond,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_iftrue,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_iffalse,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094 : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_return_output);

-- rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_cond,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_iftrue,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_iffalse,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396 : entity work.BIN_OP_EQ_uint3_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_return_output);

-- rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_cond,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_iftrue,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_iffalse,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 elem_val,
 ref_toks_0,
 var_dim_0,
 -- All submodule outputs
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_return_output,
 rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_return_output,
 rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_return_output,
 rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_return_output,
 rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_return_output,
 rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_return_output,
 rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_return_output,
 rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_return_output,
 rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_elem_val : unsigned(7 downto 0);
 variable VAR_ref_toks_0 : uint8_t_8;
 variable VAR_var_dim_0 : unsigned(2 downto 0);
 variable VAR_return_output : uint8_t_array_8_t;
 variable VAR_base : uint8_t_8;
 variable VAR_rv : uint8_t_array_8_t;
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_2c5c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_a68e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_6721_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_1b7c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_3e6b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_ef06_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_eaa4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_346f_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_e759_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_8d9c_return_output : uint8_t_array_8_t;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_elem_val := elem_val;
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_iftrue := VAR_elem_val;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_iftrue := VAR_elem_val;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_iftrue := VAR_elem_val;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_iftrue := VAR_elem_val;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_iftrue := VAR_elem_val;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_iftrue := VAR_elem_val;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_iftrue := VAR_elem_val;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_iftrue := VAR_elem_val;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_left := VAR_var_dim_0;
     -- CONST_REF_RD_uint8_t_uint8_t_8_7_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_3e6b] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_3e6b_return_output := VAR_ref_toks_0(7);

     -- CONST_REF_RD_uint8_t_uint8_t_8_4_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_1b7c] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_1b7c_return_output := VAR_ref_toks_0(4);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_2_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_2c5c] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_2c5c_return_output := VAR_ref_toks_0(2);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_0_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_ef06] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_ef06_return_output := VAR_ref_toks_0(0);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_6_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_eaa4] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_eaa4_return_output := VAR_ref_toks_0(6);

     -- CONST_REF_RD_uint8_t_uint8_t_8_3_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_346f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_346f_return_output := VAR_ref_toks_0(3);

     -- CONST_REF_RD_uint8_t_uint8_t_8_1_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_6721] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_6721_return_output := VAR_ref_toks_0(1);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_5_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_a68e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_a68e_return_output := VAR_ref_toks_0(5);

     -- Submodule level 1
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_3ec8_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_73ef_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_0c15_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_700f_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_fcd7_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_0a46_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_4094_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_c396_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_ef06_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_6721_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_2c5c_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_346f_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_1b7c_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_a68e_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_eaa4_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_3e6b_return_output;
     -- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678] LATENCY=0
     -- Inputs
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_cond <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_cond;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_iftrue <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_iftrue;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_iffalse <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_iffalse;
     -- Outputs
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_return_output := rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_return_output;

     -- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531] LATENCY=0
     -- Inputs
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_cond <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_cond;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_iftrue <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_iftrue;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_iffalse <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_iffalse;
     -- Outputs
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_return_output := rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_return_output;

     -- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea] LATENCY=0
     -- Inputs
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_cond <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_cond;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_iftrue <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_iftrue;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_iffalse <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_iffalse;
     -- Outputs
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_return_output := rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_return_output;

     -- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412] LATENCY=0
     -- Inputs
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_cond <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_cond;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_iftrue <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_iftrue;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_iffalse <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_iffalse;
     -- Outputs
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_return_output := rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_return_output;

     -- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913] LATENCY=0
     -- Inputs
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_cond <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_cond;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_iftrue <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_iftrue;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_iffalse <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_iffalse;
     -- Outputs
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_return_output := rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_return_output;

     -- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a] LATENCY=0
     -- Inputs
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_cond <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_cond;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_iftrue <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_iftrue;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_iffalse <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_iffalse;
     -- Outputs
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_return_output := rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_return_output;

     -- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43] LATENCY=0
     -- Inputs
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_cond <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_cond;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_iftrue <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_iftrue;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_iffalse <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_iffalse;
     -- Outputs
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_return_output := rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_return_output;

     -- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859] LATENCY=0
     -- Inputs
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_cond <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_cond;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_iftrue <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_iftrue;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_iffalse <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_iffalse;
     -- Outputs
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_return_output := rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_return_output;

     -- Submodule level 2
     -- CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_e759[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_8d9c] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_e759_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_8d9c_return_output := CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_e759(
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_ca43_return_output,
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_3bea_return_output,
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d913_return_output,
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_3412_return_output,
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_7859_return_output,
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_d63a_return_output,
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_8678_return_output,
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_2531_return_output);

     -- Submodule level 3
     VAR_return_output := VAR_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_e759_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_8d9c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
