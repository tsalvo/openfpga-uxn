-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 43
entity opc_div_phased_0CLK_64632f92 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_div_phased_0CLK_64632f92;
architecture arch of opc_div_phased_0CLK_64632f92 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l1101_c6_f727]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1101_c1_bf88]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1104_c7_ae9e]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1101_c2_6835]
signal t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1101_c2_6835]
signal n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1101_c2_6835]
signal result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output : unsigned(0 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l1102_c12_2632]
signal set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1104_c11_6695]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1104_c1_9d0f]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1107_c7_298b]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1104_c7_ae9e]
signal t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1104_c7_ae9e]
signal n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1104_c7_ae9e]
signal result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output : unsigned(0 downto 0);

-- t_register[uxn_opcodes_phased_h_l1105_c8_7cd6]
signal t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_stack_ptr : unsigned(7 downto 0);
signal t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1107_c11_89d1]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1107_c1_0d9d]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1110_c7_1975]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1107_c7_298b]
signal t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1107_c7_298b]
signal n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1107_c7_298b]
signal result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l1108_c8_9c84]
signal n_register_uxn_opcodes_phased_h_l1108_c8_9c84_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1108_c8_9c84_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1108_c8_9c84_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l1108_c8_9c84_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1110_c11_a9a6]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1110_c1_c298]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1113_c7_b42d]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1110_c7_1975]
signal n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1110_c7_1975]
signal result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l1111_c8_396f]
signal n_register_uxn_opcodes_phased_h_l1111_c8_396f_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1111_c8_396f_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1111_c8_396f_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l1111_c8_396f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1113_c11_557d]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1113_c1_c162]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1116_c7_e2d5]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1113_c7_b42d]
signal result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output : unsigned(0 downto 0);

-- set[uxn_opcodes_phased_h_l1114_c3_8e34]
signal set_uxn_opcodes_phased_h_l1114_c3_8e34_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l1114_c3_8e34_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1114_c3_8e34_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l1114_c3_8e34_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1114_c3_8e34_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1114_c3_8e34_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1114_c3_8e34_add : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1116_c11_0072]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1119_c7_7b91]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1116_c7_e2d5]
signal result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1117_c12_ab0c]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1119_c11_1a23]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1119_c1_3c6c]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1119_c7_7b91]
signal result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output : unsigned(0 downto 0);

-- BIN_OP_DIV[uxn_opcodes_phased_h_l1120_c33_f4bd]
signal BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_left : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_right : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_return_output : unsigned(7 downto 0);

-- put_stack[uxn_opcodes_phased_h_l1120_c3_c941]
signal put_stack_uxn_opcodes_phased_h_l1120_c3_c941_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1120_c3_c941_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1120_c3_c941_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1120_c3_c941_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1120_c3_c941_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1122_c11_2a0c]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1122_c7_2450]
signal result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727
BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835
t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond,
t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835
n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond,
n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1101_c2_6835
result_MUX_uxn_opcodes_phased_h_l1101_c2_6835 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond,
result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue,
result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse,
result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632
set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632 : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_sp,
set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_k,
set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_mul,
set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_add,
set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695
BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e
t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond,
t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e
n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond,
n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e
result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond,
result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue,
result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse,
result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output);

-- t_register_uxn_opcodes_phased_h_l1105_c8_7cd6
t_register_uxn_opcodes_phased_h_l1105_c8_7cd6 : entity work.t_register_0CLK_621d5f60 port map (
clk,
t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_CLOCK_ENABLE,
t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_stack_index,
t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_stack_ptr,
t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1
BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b
t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond,
t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b
n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond,
n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1107_c7_298b
result_MUX_uxn_opcodes_phased_h_l1107_c7_298b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond,
result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue,
result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse,
result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output);

-- n_register_uxn_opcodes_phased_h_l1108_c8_9c84
n_register_uxn_opcodes_phased_h_l1108_c8_9c84 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l1108_c8_9c84_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l1108_c8_9c84_stack_index,
n_register_uxn_opcodes_phased_h_l1108_c8_9c84_stack_ptr,
n_register_uxn_opcodes_phased_h_l1108_c8_9c84_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6
BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975
n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond,
n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1110_c7_1975
result_MUX_uxn_opcodes_phased_h_l1110_c7_1975 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond,
result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue,
result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse,
result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output);

-- n_register_uxn_opcodes_phased_h_l1111_c8_396f
n_register_uxn_opcodes_phased_h_l1111_c8_396f : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l1111_c8_396f_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l1111_c8_396f_stack_index,
n_register_uxn_opcodes_phased_h_l1111_c8_396f_stack_ptr,
n_register_uxn_opcodes_phased_h_l1111_c8_396f_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d
BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d
result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_cond,
result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iftrue,
result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iffalse,
result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output);

-- set_uxn_opcodes_phased_h_l1114_c3_8e34
set_uxn_opcodes_phased_h_l1114_c3_8e34 : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l1114_c3_8e34_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l1114_c3_8e34_sp,
set_uxn_opcodes_phased_h_l1114_c3_8e34_stack_index,
set_uxn_opcodes_phased_h_l1114_c3_8e34_ins,
set_uxn_opcodes_phased_h_l1114_c3_8e34_k,
set_uxn_opcodes_phased_h_l1114_c3_8e34_mul,
set_uxn_opcodes_phased_h_l1114_c3_8e34_add);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072
BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5
result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_cond,
result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iftrue,
result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iffalse,
result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c
BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23
BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91
result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_cond,
result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iftrue,
result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iffalse,
result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output);

-- BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd
BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd : entity work.BIN_OP_DIV_uint8_t_uint8_t_0CLK_a148083c port map (
BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_left,
BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_right,
BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_return_output);

-- put_stack_uxn_opcodes_phased_h_l1120_c3_c941
put_stack_uxn_opcodes_phased_h_l1120_c3_c941 : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l1120_c3_c941_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l1120_c3_c941_sp,
put_stack_uxn_opcodes_phased_h_l1120_c3_c941_stack_index,
put_stack_uxn_opcodes_phased_h_l1120_c3_c941_offset,
put_stack_uxn_opcodes_phased_h_l1120_c3_c941_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c
BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1122_c7_2450
result_MUX_uxn_opcodes_phased_h_l1122_c7_2450 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_cond,
result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_iftrue,
result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_iffalse,
result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 n8,
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output,
 result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output,
 set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output,
 result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output,
 t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output,
 result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output,
 n_register_uxn_opcodes_phased_h_l1108_c8_9c84_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output,
 result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output,
 n_register_uxn_opcodes_phased_h_l1111_c8_396f_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output,
 result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output,
 result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_return_output,
 result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output,
 BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_return_output,
 result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_stack_ptr : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1108_c8_9c84_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1108_c8_9c84_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1108_c8_9c84_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1108_c8_9c84_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1111_c8_396f_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1111_c8_396f_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1111_c8_396f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1111_c8_396f_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_cond : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_value : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_return_output : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_n8 := n8;
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_offset := resize(to_unsigned(0, 1), 8);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_right := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_add := resize(to_signed(-1, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_right := to_unsigned(2, 2);
     VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_mul := resize(to_unsigned(2, 2), 8);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_iffalse := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_mul := resize(to_unsigned(2, 2), 8);
     VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_add := resize(to_signed(-1, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_right := to_unsigned(5, 3);
     VAR_result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_right := to_unsigned(3, 2);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_right := to_unsigned(4, 3);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_iffalse := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_iffalse := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_k := VAR_k;
     VAR_BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_left := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_left := VAR_phase;
     VAR_result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_iffalse := result;
     VAR_n_register_uxn_opcodes_phased_h_l1108_c8_9c84_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l1111_c8_396f_stack_ptr := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_sp := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_sp := VAR_sp;
     VAR_t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l1108_c8_9c84_stack_index := VAR_stack_index;
     VAR_n_register_uxn_opcodes_phased_h_l1111_c8_396f_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_stack_index := VAR_stack_index;
     VAR_BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_right := t8;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_left := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1117_c12_ab0c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1122_c11_2a0c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1116_c11_0072] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1113_c11_557d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1110_c11_a9a6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1104_c11_6695] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1119_c11_1a23] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1107_c11_89d1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_return_output;

     -- BIN_OP_DIV[uxn_opcodes_phased_h_l1120_c33_f4bd] LATENCY=0
     -- Inputs
     BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_left <= VAR_BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_left;
     BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_right <= VAR_BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_right;
     -- Outputs
     VAR_BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_return_output := BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1101_c6_f727] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_return_output;

     -- Submodule level 1
     VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_value := VAR_BIN_OP_DIV_uxn_opcodes_phased_h_l1120_c33_f4bd_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1101_c6_f727_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1104_c11_6695_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1107_c11_89d1_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1110_c11_a9a6_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1113_c11_557d_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1116_c11_0072_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iftrue := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1117_c12_ab0c_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1119_c11_1a23_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1122_c11_2a0c_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1104_c7_ae9e] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1101_c1_bf88] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1122_c7_2450] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_cond;
     result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_return_output := result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1101_c1_bf88_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1122_c7_2450_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1107_c7_298b] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1104_c1_9d0f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_return_output;

     -- set_will_fail[uxn_opcodes_phased_h_l1102_c12_2632] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_sp;
     set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_k;
     set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_mul;
     set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_return_output := set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1119_c7_7b91] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_cond;
     result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output := result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output;
     VAR_t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1104_c1_9d0f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l1102_c12_2632_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l1116_c7_e2d5] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_cond;
     result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output := result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1110_c7_1975] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output;

     -- t_register[uxn_opcodes_phased_h_l1105_c8_7cd6] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_stack_index <= VAR_t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_stack_index;
     t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_stack_ptr <= VAR_t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_stack_ptr;
     -- Outputs
     VAR_t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_return_output := t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1107_c1_0d9d] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l1108_c8_9c84_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1107_c1_0d9d_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue := VAR_t_register_uxn_opcodes_phased_h_l1105_c8_7cd6_return_output;
     -- n_register[uxn_opcodes_phased_h_l1108_c8_9c84] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l1108_c8_9c84_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l1108_c8_9c84_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l1108_c8_9c84_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l1108_c8_9c84_stack_index;
     n_register_uxn_opcodes_phased_h_l1108_c8_9c84_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l1108_c8_9c84_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l1108_c8_9c84_return_output := n_register_uxn_opcodes_phased_h_l1108_c8_9c84_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1113_c7_b42d] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1113_c7_b42d] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_cond;
     result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output := result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1110_c1_c298] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_return_output;

     -- Submodule level 5
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l1111_c8_396f_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1110_c1_c298_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue := VAR_n_register_uxn_opcodes_phased_h_l1108_c8_9c84_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1113_c7_b42d_return_output;
     -- n_register[uxn_opcodes_phased_h_l1111_c8_396f] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l1111_c8_396f_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l1111_c8_396f_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l1111_c8_396f_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l1111_c8_396f_stack_index;
     n_register_uxn_opcodes_phased_h_l1111_c8_396f_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l1111_c8_396f_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l1111_c8_396f_return_output := n_register_uxn_opcodes_phased_h_l1111_c8_396f_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1110_c7_1975] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond;
     result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output := result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1116_c7_e2d5] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1113_c1_c162] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l1107_c7_298b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond;
     t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output := t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output;

     -- Submodule level 6
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1116_c7_e2d5_return_output;
     VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1113_c1_c162_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue := VAR_n_register_uxn_opcodes_phased_h_l1111_c8_396f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output;
     -- t8_MUX[uxn_opcodes_phased_h_l1104_c7_ae9e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond;
     t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output := t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1107_c7_298b] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond;
     result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output := result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output;

     -- set[uxn_opcodes_phased_h_l1114_c3_8e34] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l1114_c3_8e34_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l1114_c3_8e34_sp <= VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_sp;
     set_uxn_opcodes_phased_h_l1114_c3_8e34_stack_index <= VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_stack_index;
     set_uxn_opcodes_phased_h_l1114_c3_8e34_ins <= VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_ins;
     set_uxn_opcodes_phased_h_l1114_c3_8e34_k <= VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_k;
     set_uxn_opcodes_phased_h_l1114_c3_8e34_mul <= VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_mul;
     set_uxn_opcodes_phased_h_l1114_c3_8e34_add <= VAR_set_uxn_opcodes_phased_h_l1114_c3_8e34_add;
     -- Outputs

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1119_c7_7b91] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output;

     -- n8_MUX[uxn_opcodes_phased_h_l1110_c7_1975] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_cond;
     n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output := n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output;

     -- Submodule level 7
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c7_7b91_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1110_c7_1975_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l1104_c7_ae9e] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond;
     result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output := result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1119_c1_3c6c] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l1101_c2_6835] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond;
     t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output := t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output;

     -- n8_MUX[uxn_opcodes_phased_h_l1107_c7_298b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_cond;
     n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output := n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output;

     -- Submodule level 8
     VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1119_c1_3c6c_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1107_c7_298b_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1104_c7_ae9e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_cond;
     n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output := n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1101_c2_6835] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond;
     result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output := result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output;

     -- put_stack[uxn_opcodes_phased_h_l1120_c3_c941] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l1120_c3_c941_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l1120_c3_c941_sp <= VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_sp;
     put_stack_uxn_opcodes_phased_h_l1120_c3_c941_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_stack_index;
     put_stack_uxn_opcodes_phased_h_l1120_c3_c941_offset <= VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_offset;
     put_stack_uxn_opcodes_phased_h_l1120_c3_c941_value <= VAR_put_stack_uxn_opcodes_phased_h_l1120_c3_c941_value;
     -- Outputs

     -- Submodule level 9
     VAR_n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1104_c7_ae9e_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1101_c2_6835] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_cond;
     n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output := n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output;

     -- Submodule level 10
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_phased_h_l1101_c2_6835_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     n8 <= REG_COMB_n8;
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
