-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity ovr_0CLK_61914e8d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ovr_0CLK_61914e8d;
architecture arch of ovr_0CLK_61914e8d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l297_c6_b6be]
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l297_c2_2ffe]
signal n8_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l297_c2_2ffe]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l297_c2_2ffe]
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l297_c2_2ffe]
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l297_c2_2ffe]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l297_c2_2ffe]
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l297_c2_2ffe]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l297_c2_2ffe]
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l297_c2_2ffe]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l297_c2_2ffe]
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l297_c2_2ffe]
signal t8_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l310_c11_a21e]
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l310_c7_e1a4]
signal n8_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l310_c7_e1a4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l310_c7_e1a4]
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l310_c7_e1a4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l310_c7_e1a4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l310_c7_e1a4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l310_c7_e1a4]
signal t8_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l313_c11_ec0c]
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l313_c7_9648]
signal n8_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_9648_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l313_c7_9648]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l313_c7_9648]
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l313_c7_9648]
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l313_c7_9648]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l313_c7_9648]
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l313_c7_9648]
signal t8_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_9648_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l315_c30_001f]
signal sp_relative_shift_uxn_opcodes_h_l315_c30_001f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_001f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_001f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_001f_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l320_c11_3a4a]
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l320_c7_7ad5]
signal n8_MUX_uxn_opcodes_h_l320_c7_7ad5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l320_c7_7ad5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l320_c7_7ad5]
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l320_c7_7ad5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l320_c7_7ad5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l326_c11_63c3]
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l326_c7_b233]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l326_c7_b233]
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l326_c7_b233]
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_b856( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be
BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_left,
BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_right,
BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output);

-- n8_MUX_uxn_opcodes_h_l297_c2_2ffe
n8_MUX_uxn_opcodes_h_l297_c2_2ffe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l297_c2_2ffe_cond,
n8_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue,
n8_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse,
n8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe
result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_cond,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output);

-- t8_MUX_uxn_opcodes_h_l297_c2_2ffe
t8_MUX_uxn_opcodes_h_l297_c2_2ffe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l297_c2_2ffe_cond,
t8_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue,
t8_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse,
t8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e
BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_left,
BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_right,
BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_return_output);

-- n8_MUX_uxn_opcodes_h_l310_c7_e1a4
n8_MUX_uxn_opcodes_h_l310_c7_e1a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l310_c7_e1a4_cond,
n8_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue,
n8_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse,
n8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4
result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_cond,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output);

-- t8_MUX_uxn_opcodes_h_l310_c7_e1a4
t8_MUX_uxn_opcodes_h_l310_c7_e1a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l310_c7_e1a4_cond,
t8_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue,
t8_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse,
t8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c
BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_left,
BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_right,
BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_return_output);

-- n8_MUX_uxn_opcodes_h_l313_c7_9648
n8_MUX_uxn_opcodes_h_l313_c7_9648 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l313_c7_9648_cond,
n8_MUX_uxn_opcodes_h_l313_c7_9648_iftrue,
n8_MUX_uxn_opcodes_h_l313_c7_9648_iffalse,
n8_MUX_uxn_opcodes_h_l313_c7_9648_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648
result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_cond,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_return_output);

-- t8_MUX_uxn_opcodes_h_l313_c7_9648
t8_MUX_uxn_opcodes_h_l313_c7_9648 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l313_c7_9648_cond,
t8_MUX_uxn_opcodes_h_l313_c7_9648_iftrue,
t8_MUX_uxn_opcodes_h_l313_c7_9648_iffalse,
t8_MUX_uxn_opcodes_h_l313_c7_9648_return_output);

-- sp_relative_shift_uxn_opcodes_h_l315_c30_001f
sp_relative_shift_uxn_opcodes_h_l315_c30_001f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l315_c30_001f_ins,
sp_relative_shift_uxn_opcodes_h_l315_c30_001f_x,
sp_relative_shift_uxn_opcodes_h_l315_c30_001f_y,
sp_relative_shift_uxn_opcodes_h_l315_c30_001f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a
BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_left,
BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_right,
BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_return_output);

-- n8_MUX_uxn_opcodes_h_l320_c7_7ad5
n8_MUX_uxn_opcodes_h_l320_c7_7ad5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l320_c7_7ad5_cond,
n8_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue,
n8_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse,
n8_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5
result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_cond,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3
BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_left,
BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_right,
BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233
result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_cond,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output,
 n8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
 t8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_return_output,
 n8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output,
 t8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_return_output,
 n8_MUX_uxn_opcodes_h_l313_c7_9648_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_return_output,
 t8_MUX_uxn_opcodes_h_l313_c7_9648_return_output,
 sp_relative_shift_uxn_opcodes_h_l315_c30_001f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_return_output,
 n8_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_b695 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_ef38 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_2ffe_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_9648_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_9f91 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_9648_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_e1a4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_afff : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_9648_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_9648_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_9648_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_001f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_001f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_001f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_001f_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_7ad5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_59d0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l321_c3_f0d2 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_9042 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_b233_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l310_l326_l297_DUPLICATE_44e7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_300c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l310_l320_DUPLICATE_c723_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_d1ce_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l332_l293_DUPLICATE_38b2_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_59d0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_59d0;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_001f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_9042 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_9042;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l321_c3_f0d2 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l321_c3_f0d2;
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_001f_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_9f91 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_9f91;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_b695 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_b695;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_ef38 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_ef38;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_afff := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_afff;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_001f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_9648_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse := n8;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_9648_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_9648_iffalse := t8;
     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_2ffe_return_output := result.is_stack_index_flipped;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_2ffe_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_d1ce LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_d1ce_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l310_l320_DUPLICATE_c723 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l310_l320_DUPLICATE_c723_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l310_l326_l297_DUPLICATE_44e7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l310_l326_l297_DUPLICATE_44e7_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l297_c6_b6be] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_left;
     BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output := BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l326_c7_b233] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_b233_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l313_c11_ec0c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_left;
     BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_return_output := BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l310_c11_a21e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_left;
     BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_return_output := BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l326_c11_63c3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_left;
     BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_return_output := BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l320_c11_3a4a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_left;
     BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_return_output := BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l315_c30_001f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l315_c30_001f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_001f_ins;
     sp_relative_shift_uxn_opcodes_h_l315_c30_001f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_001f_x;
     sp_relative_shift_uxn_opcodes_h_l315_c30_001f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_001f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_001f_return_output := sp_relative_shift_uxn_opcodes_h_l315_c30_001f_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_2ffe_return_output := result.is_vram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_2ffe_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_300c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_300c_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_2ffe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_2ffe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_b6be_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_e1a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_e1a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_a21e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_9648_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_9648_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_ec0c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_7ad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_3a4a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_63c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l310_l320_DUPLICATE_c723_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l310_l320_DUPLICATE_c723_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_d1ce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_d1ce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_d1ce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l310_l326_l313_l320_DUPLICATE_d1ce_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_300c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_300c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l310_l326_l297_DUPLICATE_44e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l310_l326_l297_DUPLICATE_44e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l310_l326_l297_DUPLICATE_44e7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_2ffe_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_2ffe_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_2ffe_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_2ffe_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_b233_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_001f_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l326_c7_b233] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output;

     -- n8_MUX[uxn_opcodes_h_l320_c7_7ad5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l320_c7_7ad5_cond <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_7ad5_cond;
     n8_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue;
     n8_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output := n8_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l326_c7_b233] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l326_c7_b233] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_cond;
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_return_output := result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l313_c7_9648] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_return_output;

     -- t8_MUX[uxn_opcodes_h_l313_c7_9648] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l313_c7_9648_cond <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_9648_cond;
     t8_MUX_uxn_opcodes_h_l313_c7_9648_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_9648_iftrue;
     t8_MUX_uxn_opcodes_h_l313_c7_9648_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_9648_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_9648_return_output := t8_MUX_uxn_opcodes_h_l313_c7_9648_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l320_c7_7ad5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_9648_iffalse := VAR_n8_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_b233_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_9648_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_b233_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_b233_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse := VAR_t8_MUX_uxn_opcodes_h_l313_c7_9648_return_output;
     -- t8_MUX[uxn_opcodes_h_l310_c7_e1a4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l310_c7_e1a4_cond <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_e1a4_cond;
     t8_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue;
     t8_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output := t8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;

     -- n8_MUX[uxn_opcodes_h_l313_c7_9648] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l313_c7_9648_cond <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_9648_cond;
     n8_MUX_uxn_opcodes_h_l313_c7_9648_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_9648_iftrue;
     n8_MUX_uxn_opcodes_h_l313_c7_9648_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_9648_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_9648_return_output := n8_MUX_uxn_opcodes_h_l313_c7_9648_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l320_c7_7ad5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l313_c7_9648] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l320_c7_7ad5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l320_c7_7ad5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output := result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l310_c7_e1a4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse := VAR_n8_MUX_uxn_opcodes_h_l313_c7_9648_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_9648_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_7ad5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse := VAR_t8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;
     -- t8_MUX[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l297_c2_2ffe_cond <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_2ffe_cond;
     t8_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue;
     t8_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output := t8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output;

     -- n8_MUX[uxn_opcodes_h_l310_c7_e1a4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l310_c7_e1a4_cond <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_e1a4_cond;
     n8_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue;
     n8_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output := n8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l310_c7_e1a4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l313_c7_9648] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_cond;
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_return_output := result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l313_c7_9648] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l313_c7_9648] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse := VAR_n8_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_9648_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_9648_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_9648_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l310_c7_e1a4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output := result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output;

     -- n8_MUX[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l297_c2_2ffe_cond <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_2ffe_cond;
     n8_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue;
     n8_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output := n8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l310_c7_e1a4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l310_c7_e1a4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_e1a4_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_cond;
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output := result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l297_c2_2ffe] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l332_l293_DUPLICATE_38b2 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l332_l293_DUPLICATE_38b2_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_b856(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_2ffe_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l332_l293_DUPLICATE_38b2_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l332_l293_DUPLICATE_38b2_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
