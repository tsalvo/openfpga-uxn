-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 48
entity swp_0CLK_faaf4b1a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end swp_0CLK_faaf4b1a;
architecture arch of swp_0CLK_faaf4b1a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2406_c6_692c]
signal BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2406_c1_b738]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2406_c2_e90e]
signal n8_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2406_c2_e90e]
signal t8_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2406_c2_e90e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2406_c2_e90e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2406_c2_e90e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2406_c2_e90e]
signal result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2406_c2_e90e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2406_c2_e90e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l2407_c3_83cd[uxn_opcodes_h_l2407_c3_83cd]
signal printf_uxn_opcodes_h_l2407_c3_83cd_uxn_opcodes_h_l2407_c3_83cd_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2411_c11_c695]
signal BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2411_c7_91ed]
signal n8_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2411_c7_91ed]
signal t8_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2411_c7_91ed]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2411_c7_91ed]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2411_c7_91ed]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2411_c7_91ed]
signal result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2411_c7_91ed]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2411_c7_91ed]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2414_c11_63df]
signal BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2414_c7_0cd8]
signal n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2414_c7_0cd8]
signal t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2414_c7_0cd8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2414_c7_0cd8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2414_c7_0cd8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2414_c7_0cd8]
signal result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2414_c7_0cd8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2414_c7_0cd8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2417_c11_aa76]
signal BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2417_c7_34b6]
signal n8_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2417_c7_34b6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2417_c7_34b6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2417_c7_34b6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2417_c7_34b6]
signal result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2417_c7_34b6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2417_c7_34b6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2420_c30_b870]
signal sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2425_c11_a68c]
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2425_c7_d4b5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2425_c7_d4b5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2425_c7_d4b5]
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2425_c7_d4b5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2425_c7_d4b5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2430_c11_e498]
signal BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2430_c7_4fe2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2430_c7_4fe2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c551( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c
BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_left,
BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_right,
BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_return_output);

-- n8_MUX_uxn_opcodes_h_l2406_c2_e90e
n8_MUX_uxn_opcodes_h_l2406_c2_e90e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2406_c2_e90e_cond,
n8_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue,
n8_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse,
n8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output);

-- t8_MUX_uxn_opcodes_h_l2406_c2_e90e
t8_MUX_uxn_opcodes_h_l2406_c2_e90e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2406_c2_e90e_cond,
t8_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue,
t8_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse,
t8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e
result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e
result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e
result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e
result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output);

-- printf_uxn_opcodes_h_l2407_c3_83cd_uxn_opcodes_h_l2407_c3_83cd
printf_uxn_opcodes_h_l2407_c3_83cd_uxn_opcodes_h_l2407_c3_83cd : entity work.printf_uxn_opcodes_h_l2407_c3_83cd_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2407_c3_83cd_uxn_opcodes_h_l2407_c3_83cd_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695
BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_left,
BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_right,
BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output);

-- n8_MUX_uxn_opcodes_h_l2411_c7_91ed
n8_MUX_uxn_opcodes_h_l2411_c7_91ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2411_c7_91ed_cond,
n8_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue,
n8_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse,
n8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output);

-- t8_MUX_uxn_opcodes_h_l2411_c7_91ed
t8_MUX_uxn_opcodes_h_l2411_c7_91ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2411_c7_91ed_cond,
t8_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue,
t8_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse,
t8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed
result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed
result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed
result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_cond,
result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed
result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed
result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df
BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_left,
BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_right,
BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output);

-- n8_MUX_uxn_opcodes_h_l2414_c7_0cd8
n8_MUX_uxn_opcodes_h_l2414_c7_0cd8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond,
n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue,
n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse,
n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output);

-- t8_MUX_uxn_opcodes_h_l2414_c7_0cd8
t8_MUX_uxn_opcodes_h_l2414_c7_0cd8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond,
t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue,
t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse,
t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8
result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8
result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8
result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8
result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76
BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_left,
BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_right,
BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_return_output);

-- n8_MUX_uxn_opcodes_h_l2417_c7_34b6
n8_MUX_uxn_opcodes_h_l2417_c7_34b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2417_c7_34b6_cond,
n8_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue,
n8_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse,
n8_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6
result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6
result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6
result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6
result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2420_c30_b870
sp_relative_shift_uxn_opcodes_h_l2420_c30_b870 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_ins,
sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_x,
sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_y,
sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c
BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_left,
BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_right,
BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond,
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498
BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_left,
BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_right,
BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2
result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2
result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_return_output,
 n8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output,
 t8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output,
 n8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output,
 t8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output,
 n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output,
 t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_return_output,
 n8_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output,
 sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2408_c3_1387 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2407_c3_83cd_uxn_opcodes_h_l2407_c3_83cd_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2412_c3_3259 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2422_c3_2f64 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2427_c3_e29b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2411_l2406_l2430_l2425_DUPLICATE_27f7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2406_l2417_l2411_l2414_DUPLICATE_6206_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_a3a6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_80f3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2417_l2414_l2411_l2430_l2425_DUPLICATE_8131_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2425_l2414_DUPLICATE_e3bf_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2435_l2402_DUPLICATE_62d4_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2408_c3_1387 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2408_c3_1387;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2427_c3_e29b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2427_c3_e29b;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2422_c3_2f64 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2422_c3_2f64;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2412_c3_3259 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2412_c3_3259;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2417_l2414_l2411_l2430_l2425_DUPLICATE_8131 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2417_l2414_l2411_l2430_l2425_DUPLICATE_8131_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_a3a6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_a3a6_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2411_c11_c695] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_left;
     BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output := BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2406_c6_692c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2414_c11_63df] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_left;
     BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output := BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2430_c11_e498] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_left;
     BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_return_output := BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2425_l2414_DUPLICATE_e3bf LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2425_l2414_DUPLICATE_e3bf_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l2420_c30_b870] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_ins;
     sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_x;
     sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_return_output := sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2425_c11_a68c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2417_c11_aa76] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_left;
     BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_return_output := BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2411_l2406_l2430_l2425_DUPLICATE_27f7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2411_l2406_l2430_l2425_DUPLICATE_27f7_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2406_l2417_l2411_l2414_DUPLICATE_6206 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2406_l2417_l2411_l2414_DUPLICATE_6206_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_80f3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_80f3_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2406_c2_e90e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2406_c2_e90e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2406_c6_692c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2411_c7_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2411_c7_91ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2411_c11_c695_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c11_63df_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2417_c7_34b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2417_c11_aa76_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_a68c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2430_c11_e498_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2406_l2417_l2411_l2414_DUPLICATE_6206_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2406_l2417_l2411_l2414_DUPLICATE_6206_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2406_l2417_l2411_l2414_DUPLICATE_6206_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2406_l2417_l2411_l2414_DUPLICATE_6206_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2417_l2414_l2411_l2430_l2425_DUPLICATE_8131_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2417_l2414_l2411_l2430_l2425_DUPLICATE_8131_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2417_l2414_l2411_l2430_l2425_DUPLICATE_8131_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2417_l2414_l2411_l2430_l2425_DUPLICATE_8131_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2417_l2414_l2411_l2430_l2425_DUPLICATE_8131_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_80f3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_80f3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_80f3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_80f3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2411_l2406_l2430_l2425_DUPLICATE_27f7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2411_l2406_l2430_l2425_DUPLICATE_27f7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2411_l2406_l2430_l2425_DUPLICATE_27f7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2411_l2406_l2430_l2425_DUPLICATE_27f7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2411_l2406_l2430_l2425_DUPLICATE_27f7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2425_l2414_DUPLICATE_e3bf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2425_l2414_DUPLICATE_e3bf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_a3a6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_a3a6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_a3a6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2406_l2411_l2425_l2414_DUPLICATE_a3a6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2420_c30_b870_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2425_c7_d4b5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output := result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2430_c7_4fe2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output;

     -- t8_MUX[uxn_opcodes_h_l2414_c7_0cd8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond <= VAR_t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond;
     t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue;
     t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output := t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2406_c1_b738] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2417_c7_34b6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2430_c7_4fe2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output;

     -- n8_MUX[uxn_opcodes_h_l2417_c7_34b6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2417_c7_34b6_cond <= VAR_n8_MUX_uxn_opcodes_h_l2417_c7_34b6_cond;
     n8_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue;
     n8_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output := n8_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2425_c7_d4b5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2425_c7_d4b5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2407_c3_83cd_uxn_opcodes_h_l2407_c3_83cd_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2406_c1_b738_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2430_c7_4fe2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;
     -- printf_uxn_opcodes_h_l2407_c3_83cd[uxn_opcodes_h_l2407_c3_83cd] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2407_c3_83cd_uxn_opcodes_h_l2407_c3_83cd_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2407_c3_83cd_uxn_opcodes_h_l2407_c3_83cd_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2417_c7_34b6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2414_c7_0cd8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2425_c7_d4b5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2417_c7_34b6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2425_c7_d4b5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output;

     -- n8_MUX[uxn_opcodes_h_l2414_c7_0cd8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond;
     n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue;
     n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output := n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;

     -- t8_MUX[uxn_opcodes_h_l2411_c7_91ed] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2411_c7_91ed_cond <= VAR_t8_MUX_uxn_opcodes_h_l2411_c7_91ed_cond;
     t8_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue;
     t8_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output := t8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2417_c7_34b6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d4b5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2414_c7_0cd8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2414_c7_0cd8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2414_c7_0cd8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2417_c7_34b6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2411_c7_91ed] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;

     -- n8_MUX[uxn_opcodes_h_l2411_c7_91ed] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2411_c7_91ed_cond <= VAR_n8_MUX_uxn_opcodes_h_l2411_c7_91ed_cond;
     n8_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue;
     n8_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output := n8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2417_c7_34b6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;

     -- t8_MUX[uxn_opcodes_h_l2406_c2_e90e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2406_c2_e90e_cond <= VAR_t8_MUX_uxn_opcodes_h_l2406_c2_e90e_cond;
     t8_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue;
     t8_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output := t8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2417_c7_34b6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2411_c7_91ed] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output := result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;

     -- n8_MUX[uxn_opcodes_h_l2406_c2_e90e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2406_c2_e90e_cond <= VAR_n8_MUX_uxn_opcodes_h_l2406_c2_e90e_cond;
     n8_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue;
     n8_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output := n8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2411_c7_91ed] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2414_c7_0cd8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2414_c7_0cd8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2406_c2_e90e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2411_c7_91ed] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c7_0cd8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2411_c7_91ed] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2406_c2_e90e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2411_c7_91ed] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2406_c2_e90e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2406_c2_e90e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2411_c7_91ed_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2406_c2_e90e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2406_c2_e90e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2435_l2402_DUPLICATE_62d4 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2435_l2402_DUPLICATE_62d4_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c551(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2406_c2_e90e_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2435_l2402_DUPLICATE_62d4_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2435_l2402_DUPLICATE_62d4_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
