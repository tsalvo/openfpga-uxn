-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity ora_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ora_0CLK_64d180f1;
architecture arch of ora_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l991_c6_e13e]
signal BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l991_c2_1df3]
signal n8_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l991_c2_1df3]
signal t8_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l991_c2_1df3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l991_c2_1df3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l991_c2_1df3]
signal result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l991_c2_1df3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l991_c2_1df3]
signal result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l991_c2_1df3]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l991_c2_1df3]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l991_c2_1df3]
signal result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l991_c2_1df3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1004_c11_5249]
signal BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1004_c7_a9c3]
signal n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1004_c7_a9c3]
signal t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1004_c7_a9c3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1004_c7_a9c3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1004_c7_a9c3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1004_c7_a9c3]
signal result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1004_c7_a9c3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1007_c11_3531]
signal BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1007_c7_e223]
signal n8_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1007_c7_e223]
signal t8_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1007_c7_e223]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1007_c7_e223]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1007_c7_e223]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1007_c7_e223]
signal result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1007_c7_e223]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1010_c11_6147]
signal BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1010_c7_471c]
signal n8_MUX_uxn_opcodes_h_l1010_c7_471c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1010_c7_471c_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1010_c7_471c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1010_c7_471c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1010_c7_471c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1010_c7_471c]
signal result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1010_c7_471c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1012_c30_e6a7]
signal sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l1015_c21_e3a7]
signal BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_left : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_right : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a6df( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_vram_write := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e
BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_left,
BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_right,
BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output);

-- n8_MUX_uxn_opcodes_h_l991_c2_1df3
n8_MUX_uxn_opcodes_h_l991_c2_1df3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l991_c2_1df3_cond,
n8_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue,
n8_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse,
n8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output);

-- t8_MUX_uxn_opcodes_h_l991_c2_1df3
t8_MUX_uxn_opcodes_h_l991_c2_1df3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l991_c2_1df3_cond,
t8_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue,
t8_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse,
t8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3
result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3
result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_cond,
result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3
result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3
result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3
result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3
result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3
result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249
BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_left,
BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_right,
BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_return_output);

-- n8_MUX_uxn_opcodes_h_l1004_c7_a9c3
n8_MUX_uxn_opcodes_h_l1004_c7_a9c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond,
n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue,
n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse,
n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output);

-- t8_MUX_uxn_opcodes_h_l1004_c7_a9c3
t8_MUX_uxn_opcodes_h_l1004_c7_a9c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond,
t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue,
t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse,
t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3
result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3
result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3
result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond,
result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3
result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531
BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_left,
BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_right,
BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_return_output);

-- n8_MUX_uxn_opcodes_h_l1007_c7_e223
n8_MUX_uxn_opcodes_h_l1007_c7_e223 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1007_c7_e223_cond,
n8_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue,
n8_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse,
n8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output);

-- t8_MUX_uxn_opcodes_h_l1007_c7_e223
t8_MUX_uxn_opcodes_h_l1007_c7_e223 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1007_c7_e223_cond,
t8_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue,
t8_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse,
t8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223
result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223
result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223
result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_cond,
result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223
result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147
BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_left,
BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_right,
BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_return_output);

-- n8_MUX_uxn_opcodes_h_l1010_c7_471c
n8_MUX_uxn_opcodes_h_l1010_c7_471c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1010_c7_471c_cond,
n8_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue,
n8_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse,
n8_MUX_uxn_opcodes_h_l1010_c7_471c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c
result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c
result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c
result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7
sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_ins,
sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_x,
sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_y,
sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7
BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7 : entity work.BIN_OP_OR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_left,
BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_right,
BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output,
 n8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
 t8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_return_output,
 n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output,
 t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_return_output,
 n8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output,
 t8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_return_output,
 n8_MUX_uxn_opcodes_h_l1010_c7_471c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_return_output,
 sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_return_output,
 BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l996_c3_aa36 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1001_c3_493b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1005_c3_082c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1010_c7_471c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1010_c7_471c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1014_c3_fcf2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l991_l1010_l1004_l1007_DUPLICATE_a1c7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_2f36_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_8865_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_13c2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1010_l1007_DUPLICATE_3384_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1019_l987_DUPLICATE_8bdb_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1014_c3_fcf2 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1014_c3_fcf2;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l996_c3_aa36 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l996_c3_aa36;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1001_c3_493b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1001_c3_493b;
     VAR_sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1005_c3_082c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1005_c3_082c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse := n8;
     VAR_n8_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse := t8;
     VAR_t8_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1010_c11_6147] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_left;
     BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_return_output := BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_8865 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_8865_return_output := result.is_opc_done;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l991_c2_1df3_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1004_c11_5249] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_left;
     BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_return_output := BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1010_l1007_DUPLICATE_3384 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1010_l1007_DUPLICATE_3384_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l991_c2_1df3_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l1012_c30_e6a7] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_ins;
     sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_x;
     sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_return_output := sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l991_l1010_l1004_l1007_DUPLICATE_a1c7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l991_l1010_l1004_l1007_DUPLICATE_a1c7_return_output := result.u8_value;

     -- BIN_OP_OR[uxn_opcodes_h_l1015_c21_e3a7] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_left;
     BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_return_output := BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l991_c2_1df3_return_output := result.is_vram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l991_c2_1df3_return_output := result.is_pc_updated;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_2f36 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_2f36_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l991_c6_e13e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_left;
     BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output := BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1007_c11_3531] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_left;
     BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_return_output := BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_13c2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_13c2_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1004_c11_5249_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1007_c7_e223_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1007_c7_e223_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1007_c11_3531_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1010_c7_471c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1010_c11_6147_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l991_c2_1df3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l991_c2_1df3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l991_c6_e13e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l1015_c21_e3a7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_2f36_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_2f36_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_2f36_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_8865_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_8865_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_8865_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_13c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_13c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1010_l1004_l1007_DUPLICATE_13c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1010_l1007_DUPLICATE_3384_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1010_l1007_DUPLICATE_3384_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l991_l1010_l1004_l1007_DUPLICATE_a1c7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l991_l1010_l1004_l1007_DUPLICATE_a1c7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l991_l1010_l1004_l1007_DUPLICATE_a1c7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l991_l1010_l1004_l1007_DUPLICATE_a1c7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l991_c2_1df3_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l991_c2_1df3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l991_c2_1df3_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l991_c2_1df3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1012_c30_e6a7_return_output;
     -- t8_MUX[uxn_opcodes_h_l1007_c7_e223] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1007_c7_e223_cond <= VAR_t8_MUX_uxn_opcodes_h_l1007_c7_e223_cond;
     t8_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue;
     t8_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output := t8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1010_c7_471c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1010_c7_471c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1010_c7_471c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1010_c7_471c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_return_output;

     -- n8_MUX[uxn_opcodes_h_l1010_c7_471c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1010_c7_471c_cond <= VAR_n8_MUX_uxn_opcodes_h_l1010_c7_471c_cond;
     n8_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue;
     n8_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1010_c7_471c_return_output := n8_MUX_uxn_opcodes_h_l1010_c7_471c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1010_c7_471c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1010_c7_471c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1010_c7_471c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1010_c7_471c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1010_c7_471c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1010_c7_471c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1010_c7_471c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1007_c7_e223] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_return_output := result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1007_c7_e223] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1007_c7_e223] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1007_c7_e223] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1007_c7_e223] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;

     -- t8_MUX[uxn_opcodes_h_l1004_c7_a9c3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond <= VAR_t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond;
     t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue;
     t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output := t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;

     -- n8_MUX[uxn_opcodes_h_l1007_c7_e223] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1007_c7_e223_cond <= VAR_n8_MUX_uxn_opcodes_h_l1007_c7_e223_cond;
     n8_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1007_c7_e223_iftrue;
     n8_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1007_c7_e223_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output := n8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1007_c7_e223_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1004_c7_a9c3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;

     -- n8_MUX[uxn_opcodes_h_l1004_c7_a9c3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond <= VAR_n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond;
     n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue;
     n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output := n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1004_c7_a9c3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1004_c7_a9c3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;

     -- t8_MUX[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l991_c2_1df3_cond <= VAR_t8_MUX_uxn_opcodes_h_l991_c2_1df3_cond;
     t8_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue;
     t8_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output := t8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1004_c7_a9c3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1004_c7_a9c3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output := result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1004_c7_a9c3_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_return_output := result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_return_output;

     -- n8_MUX[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l991_c2_1df3_cond <= VAR_n8_MUX_uxn_opcodes_h_l991_c2_1df3_cond;
     n8_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue;
     n8_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output := n8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l991_c2_1df3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l991_c2_1df3_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1019_l987_DUPLICATE_8bdb LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1019_l987_DUPLICATE_8bdb_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a6df(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l991_c2_1df3_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1019_l987_DUPLICATE_8bdb_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1019_l987_DUPLICATE_8bdb_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
