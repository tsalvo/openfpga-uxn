-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 43
entity opc_swp_phased_0CLK_8e24d567 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_swp_phased_0CLK_8e24d567;
architecture arch of opc_swp_phased_0CLK_8e24d567 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l238_c6_f61e]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l238_c1_0746]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l241_c7_e763]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l238_c2_b7ad]
signal t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l238_c2_b7ad]
signal n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l238_c2_b7ad]
signal result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output : unsigned(0 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l239_c12_28cf]
signal set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l241_c11_a049]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l241_c1_9cca]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l244_c7_43b0]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l241_c7_e763]
signal t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l241_c7_e763]
signal n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l241_c7_e763]
signal result_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output : unsigned(0 downto 0);

-- t_register[uxn_opcodes_phased_h_l242_c8_0d5d]
signal t_register_uxn_opcodes_phased_h_l242_c8_0d5d_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l242_c8_0d5d_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l242_c8_0d5d_stack_ptr : unsigned(7 downto 0);
signal t_register_uxn_opcodes_phased_h_l242_c8_0d5d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l244_c11_ddb3]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l244_c1_6e61]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l247_c7_61cb]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l244_c7_43b0]
signal t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l244_c7_43b0]
signal n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l244_c7_43b0]
signal result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l245_c8_05e3]
signal n_register_uxn_opcodes_phased_h_l245_c8_05e3_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l245_c8_05e3_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l245_c8_05e3_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l245_c8_05e3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l247_c11_c9c1]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l247_c1_0b7c]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l250_c7_a9d3]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l247_c7_61cb]
signal n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l247_c7_61cb]
signal result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l248_c8_daa0]
signal n_register_uxn_opcodes_phased_h_l248_c8_daa0_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l248_c8_daa0_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l248_c8_daa0_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l248_c8_daa0_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l250_c11_f728]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l250_c1_3da5]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l253_c7_86d3]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l250_c7_a9d3]
signal result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output : unsigned(0 downto 0);

-- set[uxn_opcodes_phased_h_l251_c3_d344]
signal set_uxn_opcodes_phased_h_l251_c3_d344_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l251_c3_d344_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l251_c3_d344_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l251_c3_d344_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l251_c3_d344_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l251_c3_d344_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l251_c3_d344_add : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l253_c11_b9a5]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l253_c1_0994]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l256_c7_8eba]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l253_c7_86d3]
signal result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output : unsigned(0 downto 0);

-- put_stack[uxn_opcodes_phased_h_l254_c3_8006]
signal put_stack_uxn_opcodes_phased_h_l254_c3_8006_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l254_c3_8006_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l254_c3_8006_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l254_c3_8006_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l254_c3_8006_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l256_c11_a491]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l256_c1_8001]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l256_c7_8eba]
signal result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output : unsigned(0 downto 0);

-- put_stack[uxn_opcodes_phased_h_l257_c3_a1f7]
signal put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l259_c11_5319]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l259_c7_c591]
signal result_MUX_uxn_opcodes_phased_h_l259_c7_c591_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l259_c7_c591_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l259_c7_c591_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l259_c7_c591_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e
BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad
t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond,
t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue,
t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse,
t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad
n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond,
n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue,
n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse,
n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output);

-- result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad
result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond,
result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue,
result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse,
result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf
set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_sp,
set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_k,
set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_mul,
set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_add,
set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049
BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l241_c7_e763
t8_MUX_uxn_opcodes_phased_h_l241_c7_e763 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond,
t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue,
t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse,
t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l241_c7_e763
n8_MUX_uxn_opcodes_phased_h_l241_c7_e763 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond,
n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue,
n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse,
n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output);

-- result_MUX_uxn_opcodes_phased_h_l241_c7_e763
result_MUX_uxn_opcodes_phased_h_l241_c7_e763 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond,
result_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue,
result_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse,
result_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output);

-- t_register_uxn_opcodes_phased_h_l242_c8_0d5d
t_register_uxn_opcodes_phased_h_l242_c8_0d5d : entity work.t_register_0CLK_621d5f60 port map (
clk,
t_register_uxn_opcodes_phased_h_l242_c8_0d5d_CLOCK_ENABLE,
t_register_uxn_opcodes_phased_h_l242_c8_0d5d_stack_index,
t_register_uxn_opcodes_phased_h_l242_c8_0d5d_stack_ptr,
t_register_uxn_opcodes_phased_h_l242_c8_0d5d_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3
BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0
t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond,
t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue,
t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse,
t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0
n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond,
n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue,
n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse,
n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output);

-- result_MUX_uxn_opcodes_phased_h_l244_c7_43b0
result_MUX_uxn_opcodes_phased_h_l244_c7_43b0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond,
result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue,
result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse,
result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output);

-- n_register_uxn_opcodes_phased_h_l245_c8_05e3
n_register_uxn_opcodes_phased_h_l245_c8_05e3 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l245_c8_05e3_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l245_c8_05e3_stack_index,
n_register_uxn_opcodes_phased_h_l245_c8_05e3_stack_ptr,
n_register_uxn_opcodes_phased_h_l245_c8_05e3_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1
BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb
n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond,
n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue,
n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse,
n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output);

-- result_MUX_uxn_opcodes_phased_h_l247_c7_61cb
result_MUX_uxn_opcodes_phased_h_l247_c7_61cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond,
result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue,
result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse,
result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output);

-- n_register_uxn_opcodes_phased_h_l248_c8_daa0
n_register_uxn_opcodes_phased_h_l248_c8_daa0 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l248_c8_daa0_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l248_c8_daa0_stack_index,
n_register_uxn_opcodes_phased_h_l248_c8_daa0_stack_ptr,
n_register_uxn_opcodes_phased_h_l248_c8_daa0_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728
BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output);

-- result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3
result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_cond,
result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iftrue,
result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iffalse,
result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output);

-- set_uxn_opcodes_phased_h_l251_c3_d344
set_uxn_opcodes_phased_h_l251_c3_d344 : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l251_c3_d344_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l251_c3_d344_sp,
set_uxn_opcodes_phased_h_l251_c3_d344_stack_index,
set_uxn_opcodes_phased_h_l251_c3_d344_ins,
set_uxn_opcodes_phased_h_l251_c3_d344_k,
set_uxn_opcodes_phased_h_l251_c3_d344_mul,
set_uxn_opcodes_phased_h_l251_c3_d344_add);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5
BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output);

-- result_MUX_uxn_opcodes_phased_h_l253_c7_86d3
result_MUX_uxn_opcodes_phased_h_l253_c7_86d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_cond,
result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iftrue,
result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iffalse,
result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output);

-- put_stack_uxn_opcodes_phased_h_l254_c3_8006
put_stack_uxn_opcodes_phased_h_l254_c3_8006 : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l254_c3_8006_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l254_c3_8006_sp,
put_stack_uxn_opcodes_phased_h_l254_c3_8006_stack_index,
put_stack_uxn_opcodes_phased_h_l254_c3_8006_offset,
put_stack_uxn_opcodes_phased_h_l254_c3_8006_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491
BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_return_output);

-- result_MUX_uxn_opcodes_phased_h_l256_c7_8eba
result_MUX_uxn_opcodes_phased_h_l256_c7_8eba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_cond,
result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iftrue,
result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iffalse,
result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output);

-- put_stack_uxn_opcodes_phased_h_l257_c3_a1f7
put_stack_uxn_opcodes_phased_h_l257_c3_a1f7 : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_sp,
put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_stack_index,
put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_offset,
put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319
BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_return_output);

-- result_MUX_uxn_opcodes_phased_h_l259_c7_c591
result_MUX_uxn_opcodes_phased_h_l259_c7_c591 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l259_c7_c591_cond,
result_MUX_uxn_opcodes_phased_h_l259_c7_c591_iftrue,
result_MUX_uxn_opcodes_phased_h_l259_c7_c591_iffalse,
result_MUX_uxn_opcodes_phased_h_l259_c7_c591_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 n8,
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output,
 t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output,
 n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output,
 result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output,
 set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output,
 t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output,
 n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output,
 result_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output,
 t_register_uxn_opcodes_phased_h_l242_c8_0d5d_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output,
 t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output,
 n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output,
 result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output,
 n_register_uxn_opcodes_phased_h_l245_c8_05e3_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output,
 n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output,
 result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output,
 n_register_uxn_opcodes_phased_h_l248_c8_daa0_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output,
 result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output,
 result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_return_output,
 result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_return_output,
 result_MUX_uxn_opcodes_phased_h_l259_c7_c591_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l242_c8_0d5d_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l242_c8_0d5d_stack_ptr : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l242_c8_0d5d_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l242_c8_0d5d_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l245_c8_05e3_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l245_c8_05e3_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l245_c8_05e3_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l245_c8_05e3_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l248_c8_daa0_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l248_c8_daa0_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l248_c8_daa0_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l248_c8_daa0_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_cond : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l251_c3_d344_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l251_c3_d344_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l251_c3_d344_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l251_c3_d344_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l251_c3_d344_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l251_c3_d344_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l251_c3_d344_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_value : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l259_c7_c591_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_value : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l259_c7_c591_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l259_c7_c591_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l259_c7_c591_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_n8 := n8;
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_right := to_unsigned(4, 3);
     VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_add := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_mul := resize(to_unsigned(2, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_right := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_right := to_unsigned(2, 2);
     VAR_set_uxn_opcodes_phased_h_l251_c3_d344_mul := resize(to_unsigned(2, 2), 8);
     VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_offset := resize(to_unsigned(1, 1), 8);
     VAR_result_MUX_uxn_opcodes_phased_h_l259_c7_c591_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_right := to_unsigned(6, 3);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_iffalse := to_unsigned(0, 1);
     VAR_set_uxn_opcodes_phased_h_l251_c3_d344_add := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_right := to_unsigned(3, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue := to_unsigned(0, 1);
     VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_offset := resize(to_unsigned(0, 1), 8);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_iffalse := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_iffalse := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_right := to_unsigned(5, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l251_c3_d344_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l251_c3_d344_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_k := VAR_k;
     VAR_n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse := n8;
     VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_value := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_left := VAR_phase;
     VAR_result_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l259_c7_c591_iffalse := result;
     VAR_n_register_uxn_opcodes_phased_h_l245_c8_05e3_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l248_c8_daa0_stack_ptr := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_sp := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_sp := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l251_c3_d344_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_sp := VAR_sp;
     VAR_t_register_uxn_opcodes_phased_h_l242_c8_0d5d_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l245_c8_05e3_stack_index := VAR_stack_index;
     VAR_n_register_uxn_opcodes_phased_h_l248_c8_daa0_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_phased_h_l251_c3_d344_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_phased_h_l242_c8_0d5d_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_value := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_phased_h_l250_c11_f728] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l247_c11_c9c1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l244_c11_ddb3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l238_c6_f61e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l256_c11_a491] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l241_c11_a049] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l253_c11_b9a5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l259_c11_5319] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l238_c6_f61e_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l241_c11_a049_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l244_c11_ddb3_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l247_c11_c9c1_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l250_c11_f728_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l253_c11_b9a5_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l256_c11_a491_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l259_c7_c591_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l259_c11_5319_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l238_c1_0746] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l241_c7_e763] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l259_c7_c591] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l259_c7_c591_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l259_c7_c591_cond;
     result_MUX_uxn_opcodes_phased_h_l259_c7_c591_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l259_c7_c591_iftrue;
     result_MUX_uxn_opcodes_phased_h_l259_c7_c591_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l259_c7_c591_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l259_c7_c591_return_output := result_MUX_uxn_opcodes_phased_h_l259_c7_c591_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l238_c1_0746_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l259_c7_c591_return_output;
     -- set_will_fail[uxn_opcodes_phased_h_l239_c12_28cf] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_sp;
     set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_k;
     set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_mul;
     set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_return_output := set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l244_c7_43b0] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l241_c1_9cca] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l256_c7_8eba] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_cond;
     result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iftrue;
     result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output := result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output;
     VAR_t_register_uxn_opcodes_phased_h_l242_c8_0d5d_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l241_c1_9cca_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l239_c12_28cf_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l253_c7_86d3] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_cond;
     result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iftrue;
     result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output := result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l247_c7_61cb] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l244_c1_6e61] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_return_output;

     -- t_register[uxn_opcodes_phased_h_l242_c8_0d5d] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_phased_h_l242_c8_0d5d_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_phased_h_l242_c8_0d5d_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_phased_h_l242_c8_0d5d_stack_index <= VAR_t_register_uxn_opcodes_phased_h_l242_c8_0d5d_stack_index;
     t_register_uxn_opcodes_phased_h_l242_c8_0d5d_stack_ptr <= VAR_t_register_uxn_opcodes_phased_h_l242_c8_0d5d_stack_ptr;
     -- Outputs
     VAR_t_register_uxn_opcodes_phased_h_l242_c8_0d5d_return_output := t_register_uxn_opcodes_phased_h_l242_c8_0d5d_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l245_c8_05e3_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l244_c1_6e61_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue := VAR_t_register_uxn_opcodes_phased_h_l242_c8_0d5d_return_output;
     -- n_register[uxn_opcodes_phased_h_l245_c8_05e3] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l245_c8_05e3_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l245_c8_05e3_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l245_c8_05e3_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l245_c8_05e3_stack_index;
     n_register_uxn_opcodes_phased_h_l245_c8_05e3_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l245_c8_05e3_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l245_c8_05e3_return_output := n_register_uxn_opcodes_phased_h_l245_c8_05e3_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l250_c7_a9d3] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_cond;
     result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iftrue;
     result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output := result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l250_c7_a9d3] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l247_c1_0b7c] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_return_output;

     -- Submodule level 5
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l248_c8_daa0_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l247_c1_0b7c_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue := VAR_n_register_uxn_opcodes_phased_h_l245_c8_05e3_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l250_c7_a9d3_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l250_c1_3da5] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l244_c7_43b0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond;
     t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output := t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output;

     -- n_register[uxn_opcodes_phased_h_l248_c8_daa0] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l248_c8_daa0_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l248_c8_daa0_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l248_c8_daa0_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l248_c8_daa0_stack_index;
     n_register_uxn_opcodes_phased_h_l248_c8_daa0_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l248_c8_daa0_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l248_c8_daa0_return_output := n_register_uxn_opcodes_phased_h_l248_c8_daa0_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l247_c7_61cb] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond;
     result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue;
     result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output := result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l253_c7_86d3] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output;

     -- Submodule level 6
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c7_86d3_return_output;
     VAR_set_uxn_opcodes_phased_h_l251_c3_d344_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l250_c1_3da5_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue := VAR_n_register_uxn_opcodes_phased_h_l248_c8_daa0_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l247_c7_61cb] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_cond;
     n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output := n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output;

     -- set[uxn_opcodes_phased_h_l251_c3_d344] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l251_c3_d344_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l251_c3_d344_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l251_c3_d344_sp <= VAR_set_uxn_opcodes_phased_h_l251_c3_d344_sp;
     set_uxn_opcodes_phased_h_l251_c3_d344_stack_index <= VAR_set_uxn_opcodes_phased_h_l251_c3_d344_stack_index;
     set_uxn_opcodes_phased_h_l251_c3_d344_ins <= VAR_set_uxn_opcodes_phased_h_l251_c3_d344_ins;
     set_uxn_opcodes_phased_h_l251_c3_d344_k <= VAR_set_uxn_opcodes_phased_h_l251_c3_d344_k;
     set_uxn_opcodes_phased_h_l251_c3_d344_mul <= VAR_set_uxn_opcodes_phased_h_l251_c3_d344_mul;
     set_uxn_opcodes_phased_h_l251_c3_d344_add <= VAR_set_uxn_opcodes_phased_h_l251_c3_d344_add;
     -- Outputs

     -- t8_MUX[uxn_opcodes_phased_h_l241_c7_e763] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond;
     t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output := t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l256_c7_8eba] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l244_c7_43b0] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond;
     result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue;
     result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output := result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l253_c1_0994] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_return_output;

     -- Submodule level 7
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c7_8eba_return_output;
     VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l253_c1_0994_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l247_c7_61cb_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output;
     -- put_stack[uxn_opcodes_phased_h_l254_c3_8006] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l254_c3_8006_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l254_c3_8006_sp <= VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_sp;
     put_stack_uxn_opcodes_phased_h_l254_c3_8006_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_stack_index;
     put_stack_uxn_opcodes_phased_h_l254_c3_8006_offset <= VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_offset;
     put_stack_uxn_opcodes_phased_h_l254_c3_8006_value <= VAR_put_stack_uxn_opcodes_phased_h_l254_c3_8006_value;
     -- Outputs

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l256_c1_8001] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_return_output;

     -- n8_MUX[uxn_opcodes_phased_h_l244_c7_43b0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_cond;
     n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output := n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l238_c2_b7ad] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond;
     t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output := t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l241_c7_e763] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond;
     result_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue;
     result_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output := result_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output;

     -- Submodule level 8
     VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l256_c1_8001_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l244_c7_43b0_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l238_c2_b7ad] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond;
     result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue;
     result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output := result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output;

     -- put_stack[uxn_opcodes_phased_h_l257_c3_a1f7] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_sp <= VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_sp;
     put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_stack_index;
     put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_offset <= VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_offset;
     put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_value <= VAR_put_stack_uxn_opcodes_phased_h_l257_c3_a1f7_value;
     -- Outputs

     -- n8_MUX[uxn_opcodes_phased_h_l241_c7_e763] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_cond;
     n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output := n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output;

     -- Submodule level 9
     VAR_n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l241_c7_e763_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l238_c2_b7ad] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_cond;
     n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output := n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output;

     -- Submodule level 10
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_phased_h_l238_c2_b7ad_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     n8 <= REG_COMB_n8;
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
