-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 55
entity lit2_0CLK_edc09f97 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lit2_0CLK_edc09f97;
architecture arch of lit2_0CLK_edc09f97 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l214_c6_dab1]
signal BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l214_c1_7a82]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l214_c2_67f9]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l214_c2_67f9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l214_c2_67f9]
signal result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l214_c2_67f9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l214_c2_67f9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l214_c2_67f9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l214_c2_67f9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l214_c2_67f9]
signal result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(7 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l214_c2_67f9]
signal tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l215_c3_b971[uxn_opcodes_h_l215_c3_b971]
signal printf_uxn_opcodes_h_l215_c3_b971_uxn_opcodes_h_l215_c3_b971_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l221_c11_4630]
signal BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l221_c7_d7cb]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l221_c7_d7cb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l221_c7_d7cb]
signal result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l221_c7_d7cb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l221_c7_d7cb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l221_c7_d7cb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l221_c7_d7cb]
signal result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(7 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l221_c7_d7cb]
signal tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l223_c22_987d]
signal BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l225_c11_9b6e]
signal BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l225_c7_a321]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l225_c7_a321]
signal result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l225_c7_a321]
signal result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l225_c7_a321]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l225_c7_a321]
signal result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l225_c7_a321]
signal result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(7 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l225_c7_a321]
signal tmp16_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l227_c3_1ec5]
signal CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l229_c11_99c4]
signal BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l229_c7_3ddc]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l229_c7_3ddc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l229_c7_3ddc]
signal result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l229_c7_3ddc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l229_c7_3ddc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l229_c7_3ddc]
signal result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(7 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l229_c7_3ddc]
signal tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l230_c3_cec3]
signal BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l232_c22_9e46]
signal BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_right : unsigned(1 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l237_c11_fc25]
signal BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l237_c7_39f8]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l237_c7_39f8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l237_c7_39f8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l237_c7_39f8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l237_c7_39f8]
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_return_output : unsigned(7 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l240_c31_71d8]
signal CONST_SR_8_uxn_opcodes_h_l240_c31_71d8_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l240_c31_71d8_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l242_c11_c726]
signal BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l242_c7_056b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l242_c7_056b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_14ff( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.u8_value := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1
BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_left,
BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_right,
BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9
result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_cond,
result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9
result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_cond,
result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output);

-- tmp16_MUX_uxn_opcodes_h_l214_c2_67f9
tmp16_MUX_uxn_opcodes_h_l214_c2_67f9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_cond,
tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue,
tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse,
tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_return_output);

-- printf_uxn_opcodes_h_l215_c3_b971_uxn_opcodes_h_l215_c3_b971
printf_uxn_opcodes_h_l215_c3_b971_uxn_opcodes_h_l215_c3_b971 : entity work.printf_uxn_opcodes_h_l215_c3_b971_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l215_c3_b971_uxn_opcodes_h_l215_c3_b971_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630
BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_left,
BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_right,
BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb
result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_cond,
result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb
result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_cond,
result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output);

-- tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb
tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_cond,
tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue,
tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse,
tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d
BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_left,
BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_right,
BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e
BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_left,
BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_right,
BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321
result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_cond,
result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321
result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_cond,
result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output);

-- tmp16_MUX_uxn_opcodes_h_l225_c7_a321
tmp16_MUX_uxn_opcodes_h_l225_c7_a321 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l225_c7_a321_cond,
tmp16_MUX_uxn_opcodes_h_l225_c7_a321_iftrue,
tmp16_MUX_uxn_opcodes_h_l225_c7_a321_iffalse,
tmp16_MUX_uxn_opcodes_h_l225_c7_a321_return_output);

-- CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5
CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5_x,
CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4
BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_left,
BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_right,
BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc
result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_cond,
result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc
result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_cond,
result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output);

-- tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc
tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_cond,
tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue,
tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse,
tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3
BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_left,
BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_right,
BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46
BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46 : entity work.BIN_OP_PLUS_uint16_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_left,
BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_right,
BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25
BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_left,
BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_right,
BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8
result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_cond,
result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_return_output);

-- CONST_SR_8_uxn_opcodes_h_l240_c31_71d8
CONST_SR_8_uxn_opcodes_h_l240_c31_71d8 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l240_c31_71d8_x,
CONST_SR_8_uxn_opcodes_h_l240_c31_71d8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726
BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_left,
BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_right,
BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 previous_ram_read,
 -- Registers
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
 tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output,
 tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output,
 tmp16_MUX_uxn_opcodes_h_l225_c7_a321_return_output,
 CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output,
 tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output,
 BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_return_output,
 CONST_SR_8_uxn_opcodes_h_l240_c31_71d8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l217_c3_c0e9 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l214_c2_67f9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l215_c3_b971_uxn_opcodes_h_l215_c3_b971_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l221_c7_d7cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l223_c3_272d : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_a321_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_a321_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_a321_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_a321_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l232_c3_550f : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l234_c3_6763 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_return_output : unsigned(16 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l235_c21_f58c_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l239_c3_3271 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_71d8_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_71d8_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l240_c21_8243_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_42c3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_7f54_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l242_l237_l225_l221_DUPLICATE_2727_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_897d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l242_l237_l229_l225_l221_DUPLICATE_bdba_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l226_l230_DUPLICATE_5529_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l229_l225_DUPLICATE_1a5a_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_14ff_uxn_opcodes_h_l247_l209_DUPLICATE_6477_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_iffalse := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l234_c3_6763 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l234_c3_6763;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l217_c3_c0e9 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l217_c3_c0e9;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l239_c3_3271 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l239_c3_3271;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_right := to_unsigned(2, 2);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_left := VAR_pc;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_left := VAR_pc;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_left := tmp16;
     VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_71d8_x := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse := tmp16;
     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l226_l230_DUPLICATE_5529 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l226_l230_DUPLICATE_5529_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_ram_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l242_c11_c726] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_left;
     BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_return_output := BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l223_c22_987d] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_left;
     BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_return_output := BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_return_output;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l214_c2_67f9] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l214_c2_67f9_return_output := result.sp_relative_shift;

     -- result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d[uxn_opcodes_h_l221_c7_d7cb] LATENCY=0
     VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l221_c7_d7cb_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l242_l237_l229_l225_l221_DUPLICATE_bdba LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l242_l237_l229_l225_l221_DUPLICATE_bdba_return_output := result.is_opc_done;

     -- CONST_SR_8[uxn_opcodes_h_l240_c31_71d8] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l240_c31_71d8_x <= VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_71d8_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_71d8_return_output := CONST_SR_8_uxn_opcodes_h_l240_c31_71d8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l221_c11_4630] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_left;
     BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output := BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l229_l225_DUPLICATE_1a5a LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l229_l225_DUPLICATE_1a5a_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_42c3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_42c3_return_output := result.is_pc_updated;

     -- BIN_OP_PLUS[uxn_opcodes_h_l232_c22_9e46] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_left;
     BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_return_output := BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_897d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_897d_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l225_c11_9b6e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_left;
     BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_return_output := BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l242_l237_l225_l221_DUPLICATE_2727 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l242_l237_l225_l221_DUPLICATE_2727_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l229_c11_99c4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_left;
     BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_return_output := BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l214_c6_dab1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_left;
     BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output := BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_7f54 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_7f54_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l237_c11_fc25] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_left;
     BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_return_output := BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_dab1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_4630_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_a321_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_9b6e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_99c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_fc25_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_c726_return_output;
     VAR_result_u16_value_uxn_opcodes_h_l223_c3_272d := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_987d_return_output, 16);
     VAR_result_u16_value_uxn_opcodes_h_l232_c3_550f := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_9e46_return_output, 16);
     VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l226_l230_DUPLICATE_5529_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l226_l230_DUPLICATE_5529_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l229_l225_DUPLICATE_1a5a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l229_l225_DUPLICATE_1a5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l242_l237_l229_l225_l221_DUPLICATE_bdba_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l242_l237_l229_l225_l221_DUPLICATE_bdba_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l242_l237_l229_l225_l221_DUPLICATE_bdba_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l242_l237_l229_l225_l221_DUPLICATE_bdba_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l242_l237_l229_l225_l221_DUPLICATE_bdba_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_42c3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_42c3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_42c3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_42c3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l242_l237_l225_l221_DUPLICATE_2727_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l242_l237_l225_l221_DUPLICATE_2727_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l242_l237_l225_l221_DUPLICATE_2727_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l242_l237_l225_l221_DUPLICATE_2727_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l242_l237_l225_l221_DUPLICATE_2727_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_7f54_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_7f54_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_7f54_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_7f54_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_897d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_897d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_897d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l237_l225_DUPLICATE_897d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse := VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l221_c7_d7cb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l214_c2_67f9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue := VAR_result_u16_value_uxn_opcodes_h_l223_c3_272d;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue := VAR_result_u16_value_uxn_opcodes_h_l232_c3_550f;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l242_c7_056b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l221_c7_d7cb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l240_c21_8243] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l240_c21_8243_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_71d8_return_output);

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l214_c2_67f9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l242_c7_056b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l237_c7_39f8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l237_c7_39f8] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l214_c1_7a82] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l229_c7_3ddc] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_cond;
     result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output := result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l230_c3_cec3] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_left;
     BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_return_output := BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l227_c3_1ec5] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5_x <= VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5_return_output := CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5_return_output;

     -- Submodule level 2
     VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l240_c21_8243_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_a321_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_1ec5_return_output;
     VAR_printf_uxn_opcodes_h_l215_c3_b971_uxn_opcodes_h_l215_c3_b971_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_7a82_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_056b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_39f8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_056b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_39f8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l237_c7_39f8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l229_c7_3ddc] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_cond;
     tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue;
     tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output := tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l235_c21_f58c] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l235_c21_f58c_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_cec3_return_output);

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l229_c7_3ddc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l237_c7_39f8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l237_c7_39f8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_return_output := result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l225_c7_a321] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_cond;
     result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output := result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l229_c7_3ddc] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;

     -- printf_uxn_opcodes_h_l215_c3_b971[uxn_opcodes_h_l215_c3_b971] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l215_c3_b971_uxn_opcodes_h_l215_c3_b971_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l215_c3_b971_uxn_opcodes_h_l215_c3_b971_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l214_c2_67f9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l235_c21_f58c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_39f8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_39f8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_39f8_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_a321_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l221_c7_d7cb] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_cond;
     result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output := result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l225_c7_a321] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l225_c7_a321_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_a321_cond;
     tmp16_MUX_uxn_opcodes_h_l225_c7_a321_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_a321_iftrue;
     tmp16_MUX_uxn_opcodes_h_l225_c7_a321_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_a321_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_a321_return_output := tmp16_MUX_uxn_opcodes_h_l225_c7_a321_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l225_c7_a321] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l229_c7_3ddc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output := result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l229_c7_3ddc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l229_c7_3ddc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l225_c7_a321] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_a321_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_a321_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_3ddc_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_a321_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l225_c7_a321] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_cond;
     result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output := result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l214_c2_67f9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output := result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l221_c7_d7cb] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l221_c7_d7cb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l225_c7_a321] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l221_c7_d7cb] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_cond;
     tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue;
     tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output := tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l225_c7_a321] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_a321_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_a321_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_a321_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l221_c7_d7cb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output := result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l221_c7_d7cb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l214_c2_67f9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l214_c2_67f9] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l221_c7_d7cb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l214_c2_67f9] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_cond;
     tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue;
     tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_return_output := tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_d7cb_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_67f9_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l214_c2_67f9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l214_c2_67f9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output := result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l214_c2_67f9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_14ff_uxn_opcodes_h_l247_l209_DUPLICATE_6477 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_14ff_uxn_opcodes_h_l247_l209_DUPLICATE_6477_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_14ff(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_67f9_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_67f9_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_14ff_uxn_opcodes_h_l247_l209_DUPLICATE_6477_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_14ff_uxn_opcodes_h_l247_l209_DUPLICATE_6477_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
