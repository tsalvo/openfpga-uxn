-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity jsr_0CLK_0cbff8de is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr_0CLK_0cbff8de;
architecture arch of jsr_0CLK_0cbff8de is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l737_c6_2588]
signal BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l737_c2_e642]
signal result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l737_c2_e642]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l737_c2_e642]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l737_c2_e642]
signal result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l737_c2_e642]
signal result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l737_c2_e642]
signal result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l737_c2_e642]
signal result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l737_c2_e642]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l737_c2_e642]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l737_c2_e642]
signal result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(15 downto 0);

-- t8_MUX[uxn_opcodes_h_l737_c2_e642]
signal t8_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l750_c11_92be]
signal BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l750_c7_9019]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l750_c7_9019]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l750_c7_9019]
signal result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l750_c7_9019]
signal result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l750_c7_9019]
signal result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l750_c7_9019]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l750_c7_9019]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l750_c7_9019]
signal result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(15 downto 0);

-- t8_MUX[uxn_opcodes_h_l750_c7_9019]
signal t8_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l752_c30_e08a]
signal sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l754_c11_ce6c]
signal BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l754_c7_aef9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l754_c7_aef9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l754_c7_aef9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l754_c7_aef9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l754_c7_aef9]
signal result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l754_c7_aef9]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l754_c7_aef9]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l754_c7_aef9]
signal result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(15 downto 0);

-- t8_MUX[uxn_opcodes_h_l754_c7_aef9]
signal t8_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l762_c11_7b12]
signal BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l762_c7_fc58]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l762_c7_fc58]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l762_c7_fc58]
signal result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l762_c7_fc58]
signal result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l762_c7_fc58]
signal result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l762_c7_fc58]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_return_output : unsigned(0 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l765_c31_5210]
signal CONST_SR_8_uxn_opcodes_h_l765_c31_5210_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l765_c31_5210_return_output : unsigned(15 downto 0);

-- u16_add_u8_as_i8[uxn_opcodes_h_l767_c22_0fa3]
signal u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_u16 : unsigned(15 downto 0);
signal u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_u8 : unsigned(7 downto 0);
signal u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_return_output : unsigned(15 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_vram_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_ram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_stack_index_flipped := ref_toks_9;
      base.u16_value := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588
BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_left,
BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_right,
BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642
result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642
result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642
result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642
result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642
result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642
result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_cond,
result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642
result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642
result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_cond,
result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output);

-- t8_MUX_uxn_opcodes_h_l737_c2_e642
t8_MUX_uxn_opcodes_h_l737_c2_e642 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l737_c2_e642_cond,
t8_MUX_uxn_opcodes_h_l737_c2_e642_iftrue,
t8_MUX_uxn_opcodes_h_l737_c2_e642_iffalse,
t8_MUX_uxn_opcodes_h_l737_c2_e642_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be
BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_left,
BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_right,
BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019
result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_cond,
result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019
result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_cond,
result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output);

-- t8_MUX_uxn_opcodes_h_l750_c7_9019
t8_MUX_uxn_opcodes_h_l750_c7_9019 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l750_c7_9019_cond,
t8_MUX_uxn_opcodes_h_l750_c7_9019_iftrue,
t8_MUX_uxn_opcodes_h_l750_c7_9019_iffalse,
t8_MUX_uxn_opcodes_h_l750_c7_9019_return_output);

-- sp_relative_shift_uxn_opcodes_h_l752_c30_e08a
sp_relative_shift_uxn_opcodes_h_l752_c30_e08a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_ins,
sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_x,
sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_y,
sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c
BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_left,
BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_right,
BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9
result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9
result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9
result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_cond,
result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9
result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_cond,
result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output);

-- t8_MUX_uxn_opcodes_h_l754_c7_aef9
t8_MUX_uxn_opcodes_h_l754_c7_aef9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l754_c7_aef9_cond,
t8_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue,
t8_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse,
t8_MUX_uxn_opcodes_h_l754_c7_aef9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12
BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_left,
BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_right,
BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58
result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58
result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58
result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_cond,
result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58
result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_cond,
result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58
result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_return_output);

-- CONST_SR_8_uxn_opcodes_h_l765_c31_5210
CONST_SR_8_uxn_opcodes_h_l765_c31_5210 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l765_c31_5210_x,
CONST_SR_8_uxn_opcodes_h_l765_c31_5210_return_output);

-- u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3
u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3 : entity work.u16_add_u8_as_i8_0CLK_e595f783 port map (
u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_u16,
u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_u8,
u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
 t8_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output,
 t8_MUX_uxn_opcodes_h_l750_c7_9019_return_output,
 sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output,
 t8_MUX_uxn_opcodes_h_l754_c7_aef9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_return_output,
 CONST_SR_8_uxn_opcodes_h_l765_c31_5210_return_output,
 u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l747_c3_f997 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l742_c3_ed42 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l737_c2_e642_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l737_c2_e642_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l750_c7_9019_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l737_c2_e642_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l737_c2_e642_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l751_c3_accb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l750_c7_9019_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l750_c7_9019_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l754_c7_aef9_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l750_c7_9019_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l759_c3_d221 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l757_c3_2cb7 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l754_c7_aef9_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l760_c21_9ac7_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l764_c3_1893 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l762_c7_fc58_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l763_c3_52dc : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l762_c7_fc58_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l765_c31_5210_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l765_c31_5210_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l765_c21_a487_return_output : unsigned(7 downto 0);
 variable VAR_u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_u16 : unsigned(15 downto 0);
 variable VAR_u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_u8 : unsigned(7 downto 0);
 variable VAR_u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l750_l762_l737_DUPLICATE_8107_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l754_l750_l762_l737_DUPLICATE_3298_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l754_l750_l762_DUPLICATE_dcfa_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l754_l750_DUPLICATE_6c5f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l754_l750_l762_DUPLICATE_8ca0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l754_l750_DUPLICATE_5d31_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l733_l771_DUPLICATE_0595_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l759_c3_d221 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l759_c3_d221;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l747_c3_f997 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l747_c3_f997;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l751_c3_accb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l751_c3_accb;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l742_c3_ed42 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l742_c3_ed42;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_right := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l757_c3_2cb7 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l757_c3_2cb7;
     VAR_sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l763_c3_52dc := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l763_c3_52dc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l764_c3_1893 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l764_c3_1893;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_ins := VAR_ins;
     VAR_CONST_SR_8_uxn_opcodes_h_l765_c31_5210_x := VAR_pc;
     VAR_u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_u16 := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l737_c2_e642_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l750_c7_9019_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse := t8;
     VAR_u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_u8 := t8;
     -- u16_add_u8_as_i8[uxn_opcodes_h_l767_c22_0fa3] LATENCY=0
     -- Inputs
     u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_u16 <= VAR_u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_u16;
     u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_u8 <= VAR_u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_u8;
     -- Outputs
     VAR_u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_return_output := u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l754_l750_l762_l737_DUPLICATE_3298 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l754_l750_l762_l737_DUPLICATE_3298_return_output := result.u16_value;

     -- sp_relative_shift[uxn_opcodes_h_l752_c30_e08a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_ins;
     sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_x;
     sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_return_output := sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l762_c7_fc58] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l762_c7_fc58_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l754_l750_DUPLICATE_6c5f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l754_l750_DUPLICATE_6c5f_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l762_c11_7b12] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_left;
     BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_return_output := BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_return_output;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l762_c7_fc58] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l762_c7_fc58_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l737_c6_2588] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_left;
     BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output := BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l737_c2_e642] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l737_c2_e642_return_output := result.is_ram_write;

     -- CONST_SR_8[uxn_opcodes_h_l765_c31_5210] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l765_c31_5210_x <= VAR_CONST_SR_8_uxn_opcodes_h_l765_c31_5210_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l765_c31_5210_return_output := CONST_SR_8_uxn_opcodes_h_l765_c31_5210_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l760_c21_9ac7] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l760_c21_9ac7_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_pc);

     -- BIN_OP_EQ[uxn_opcodes_h_l750_c11_92be] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_left;
     BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output := BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l754_l750_DUPLICATE_5d31 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l754_l750_DUPLICATE_5d31_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l754_c11_ce6c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_left;
     BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output := BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l750_l762_l737_DUPLICATE_8107 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l750_l762_l737_DUPLICATE_8107_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l754_l750_l762_DUPLICATE_dcfa LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l754_l750_l762_DUPLICATE_dcfa_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l754_l750_l762_DUPLICATE_8ca0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l754_l750_l762_DUPLICATE_8ca0_return_output := result.is_pc_updated;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l737_c2_e642] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l737_c2_e642_return_output := result.is_vram_write;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l737_c2_e642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l737_c6_2588_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l750_c7_9019_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_92be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l754_c7_aef9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c11_ce6c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_7b12_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l760_c21_9ac7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l754_l750_l762_l737_DUPLICATE_3298_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l754_l750_l762_l737_DUPLICATE_3298_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l754_l750_l762_l737_DUPLICATE_3298_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l754_l750_l762_l737_DUPLICATE_3298_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l754_l750_l762_DUPLICATE_dcfa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l754_l750_l762_DUPLICATE_dcfa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l754_l750_l762_DUPLICATE_dcfa_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l754_l750_l762_DUPLICATE_8ca0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l754_l750_l762_DUPLICATE_8ca0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l754_l750_l762_DUPLICATE_8ca0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l754_l750_DUPLICATE_5d31_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l754_l750_DUPLICATE_5d31_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l754_l750_DUPLICATE_6c5f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l754_l750_DUPLICATE_6c5f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l750_l762_l737_DUPLICATE_8107_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l750_l762_l737_DUPLICATE_8107_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l750_l762_l737_DUPLICATE_8107_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l737_c2_e642_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l737_c2_e642_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l762_c7_fc58_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l762_c7_fc58_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l752_c30_e08a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue := VAR_u16_add_u8_as_i8_uxn_opcodes_h_l767_c22_0fa3_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l762_c7_fc58] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_cond;
     result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output := result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l762_c7_fc58] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l754_c7_aef9] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l737_c2_e642] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l754_c7_aef9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l737_c2_e642] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l762_c7_fc58] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_return_output;

     -- t8_MUX[uxn_opcodes_h_l754_c7_aef9] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l754_c7_aef9_cond <= VAR_t8_MUX_uxn_opcodes_h_l754_c7_aef9_cond;
     t8_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue;
     t8_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l754_c7_aef9_return_output := t8_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l762_c7_fc58] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l762_c7_fc58] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l765_c21_a487] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l765_c21_a487_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l765_c31_5210_return_output);

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l765_c21_a487_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_fc58_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_fc58_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_fc58_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_fc58_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l750_c7_9019_iffalse := VAR_t8_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l754_c7_aef9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l754_c7_aef9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output := result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l754_c7_aef9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;

     -- t8_MUX[uxn_opcodes_h_l750_c7_9019] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l750_c7_9019_cond <= VAR_t8_MUX_uxn_opcodes_h_l750_c7_9019_cond;
     t8_MUX_uxn_opcodes_h_l750_c7_9019_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l750_c7_9019_iftrue;
     t8_MUX_uxn_opcodes_h_l750_c7_9019_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l750_c7_9019_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l750_c7_9019_return_output := t8_MUX_uxn_opcodes_h_l750_c7_9019_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l762_c7_fc58] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_cond;
     result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output := result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l750_c7_9019] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l754_c7_aef9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l754_c7_aef9] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l750_c7_9019] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_9019_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_9019_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_fc58_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l737_c2_e642_iffalse := VAR_t8_MUX_uxn_opcodes_h_l750_c7_9019_return_output;
     -- t8_MUX[uxn_opcodes_h_l737_c2_e642] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l737_c2_e642_cond <= VAR_t8_MUX_uxn_opcodes_h_l737_c2_e642_cond;
     t8_MUX_uxn_opcodes_h_l737_c2_e642_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l737_c2_e642_iftrue;
     t8_MUX_uxn_opcodes_h_l737_c2_e642_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l737_c2_e642_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l737_c2_e642_return_output := t8_MUX_uxn_opcodes_h_l737_c2_e642_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l737_c2_e642] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l737_c2_e642] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l750_c7_9019] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_cond;
     result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output := result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l750_c7_9019] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l750_c7_9019] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l754_c7_aef9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output := result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l750_c7_9019] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l750_c7_9019] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_9019_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_9019_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_9019_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_9019_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c7_aef9_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l737_c2_e642_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l750_c7_9019] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_cond;
     result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output := result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l737_c2_e642] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l737_c2_e642] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l737_c2_e642] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_cond;
     result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output := result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l737_c2_e642] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l737_c2_e642] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_return_output;

     -- Submodule level 5
     VAR_result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_9019_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l737_c2_e642] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_cond;
     result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output := result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l733_l771_DUPLICATE_0595 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l733_l771_DUPLICATE_0595_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d(
     result,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l737_c2_e642_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l737_c2_e642_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l733_l771_DUPLICATE_0595_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dd3d_uxn_opcodes_h_l733_l771_DUPLICATE_0595_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
