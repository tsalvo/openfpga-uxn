-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 56
entity inc2_0CLK_a6885b22 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc2_0CLK_a6885b22;
architecture arch of inc2_0CLK_a6885b22 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1291_c6_b69f]
signal BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1291_c1_6d0b]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1291_c2_f936]
signal tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1291_c2_f936]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1291_c2_f936]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1291_c2_f936]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1291_c2_f936]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1291_c2_f936]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1291_c2_f936]
signal result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l1291_c2_f936]
signal t16_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l1292_c3_5656[uxn_opcodes_h_l1292_c3_5656]
signal printf_uxn_opcodes_h_l1292_c3_5656_uxn_opcodes_h_l1292_c3_5656_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1296_c11_46d4]
signal BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1296_c7_c406]
signal tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1296_c7_c406]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1296_c7_c406]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1296_c7_c406]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1296_c7_c406]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1296_c7_c406]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1296_c7_c406]
signal result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l1296_c7_c406]
signal t16_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1299_c11_0719]
signal BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1299_c7_0cc4]
signal tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1299_c7_0cc4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1299_c7_0cc4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1299_c7_0cc4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1299_c7_0cc4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1299_c7_0cc4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1299_c7_0cc4]
signal result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l1299_c7_0cc4]
signal t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l1301_c3_eebc]
signal CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1303_c11_4403]
signal BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1303_c7_4f8c]
signal tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1303_c7_4f8c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1303_c7_4f8c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1303_c7_4f8c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1303_c7_4f8c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1303_c7_4f8c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1303_c7_4f8c]
signal result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l1303_c7_4f8c]
signal t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l1304_c3_62bd]
signal BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1305_c11_9b82]
signal BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_return_output : unsigned(16 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1307_c30_c1ae]
signal sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1312_c11_6062]
signal BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1312_c7_755d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1312_c7_755d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1312_c7_755d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1312_c7_755d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1312_c7_755d]
signal result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_return_output : unsigned(7 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l1315_c31_5358]
signal CONST_SR_8_uxn_opcodes_h_l1315_c31_5358_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l1315_c31_5358_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1317_c11_1342]
signal BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1317_c7_cdaf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1317_c7_cdaf]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_8c29( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f
BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_left,
BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_right,
BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1291_c2_f936
tmp16_MUX_uxn_opcodes_h_l1291_c2_f936 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_cond,
tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue,
tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse,
tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936
result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936
result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936
result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936
result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936
result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_cond,
result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_return_output);

-- t16_MUX_uxn_opcodes_h_l1291_c2_f936
t16_MUX_uxn_opcodes_h_l1291_c2_f936 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1291_c2_f936_cond,
t16_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue,
t16_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse,
t16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output);

-- printf_uxn_opcodes_h_l1292_c3_5656_uxn_opcodes_h_l1292_c3_5656
printf_uxn_opcodes_h_l1292_c3_5656_uxn_opcodes_h_l1292_c3_5656 : entity work.printf_uxn_opcodes_h_l1292_c3_5656_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1292_c3_5656_uxn_opcodes_h_l1292_c3_5656_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4
BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_left,
BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_right,
BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1296_c7_c406
tmp16_MUX_uxn_opcodes_h_l1296_c7_c406 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_cond,
tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue,
tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse,
tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406
result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406
result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406
result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406
result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406
result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_cond,
result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_return_output);

-- t16_MUX_uxn_opcodes_h_l1296_c7_c406
t16_MUX_uxn_opcodes_h_l1296_c7_c406 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1296_c7_c406_cond,
t16_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue,
t16_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse,
t16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719
BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_left,
BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_right,
BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4
tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond,
tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue,
tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse,
tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4
result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output);

-- t16_MUX_uxn_opcodes_h_l1299_c7_0cc4
t16_MUX_uxn_opcodes_h_l1299_c7_0cc4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond,
t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue,
t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse,
t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output);

-- CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc
CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc_x,
CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403
BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_left,
BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_right,
BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c
tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond,
tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue,
tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse,
tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c
result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c
result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c
result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c
result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output);

-- t16_MUX_uxn_opcodes_h_l1303_c7_4f8c
t16_MUX_uxn_opcodes_h_l1303_c7_4f8c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond,
t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue,
t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse,
t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd
BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_left,
BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_right,
BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82
BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82 : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_left,
BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_right,
BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae
sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_ins,
sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_x,
sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_y,
sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062
BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_left,
BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_right,
BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d
result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d
result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d
result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d
result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_return_output);

-- CONST_SR_8_uxn_opcodes_h_l1315_c31_5358
CONST_SR_8_uxn_opcodes_h_l1315_c31_5358 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l1315_c31_5358_x,
CONST_SR_8_uxn_opcodes_h_l1315_c31_5358_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342
BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_left,
BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_right,
BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_return_output,
 tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_return_output,
 t16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output,
 tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_return_output,
 t16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output,
 tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output,
 t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output,
 CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output,
 tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output,
 t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output,
 BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_return_output,
 sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_return_output,
 CONST_SR_8_uxn_opcodes_h_l1315_c31_5358_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_iffalse : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1293_c3_01a6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1291_c2_f936_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1292_c3_5656_uxn_opcodes_h_l1292_c3_5656_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1297_c3_9044 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1296_c7_c406_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_uxn_opcodes_h_l1305_c3_7ebe : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1309_c3_2b69 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_return_output : unsigned(16 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1310_c21_2ef9_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1314_c3_898f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l1315_c31_5358_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l1315_c31_5358_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1315_c21_ce1e_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_1730_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1299_l1296_l1291_l1317_l1312_DUPLICATE_9bdc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1291_l1303_l1296_l1299_DUPLICATE_8b2f_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_29dc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1303_l1299_l1296_l1317_l1312_DUPLICATE_f522_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1300_l1304_DUPLICATE_a97b_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1312_l1299_DUPLICATE_00f9_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1322_l1287_DUPLICATE_4025_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1314_c3_898f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1314_c3_898f;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1309_c3_2b69 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1309_c3_2b69;
     VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1293_c3_01a6 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1293_c3_01a6;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1297_c3_9044 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1297_c3_9044;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse := t16;
     VAR_CONST_SR_8_uxn_opcodes_h_l1315_c31_5358_x := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse := tmp16;
     -- CONST_SR_8[uxn_opcodes_h_l1315_c31_5358] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l1315_c31_5358_x <= VAR_CONST_SR_8_uxn_opcodes_h_l1315_c31_5358_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l1315_c31_5358_return_output := CONST_SR_8_uxn_opcodes_h_l1315_c31_5358_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_1730 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_1730_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1296_c11_46d4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1303_l1299_l1296_l1317_l1312_DUPLICATE_f522 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1303_l1299_l1296_l1317_l1312_DUPLICATE_f522_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1303_c11_4403] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_left;
     BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output := BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1300_l1304_DUPLICATE_a97b LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1300_l1304_DUPLICATE_a97b_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- sp_relative_shift[uxn_opcodes_h_l1307_c30_c1ae] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_ins;
     sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_x;
     sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_return_output := sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_29dc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_29dc_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1291_c6_b69f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1291_l1303_l1296_l1299_DUPLICATE_8b2f LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1291_l1303_l1296_l1299_DUPLICATE_8b2f_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1299_c11_0719] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_left;
     BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output := BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1317_c11_1342] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_left;
     BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_return_output := BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1299_l1296_l1291_l1317_l1312_DUPLICATE_9bdc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1299_l1296_l1291_l1317_l1312_DUPLICATE_9bdc_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1312_l1299_DUPLICATE_00f9 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1312_l1299_DUPLICATE_00f9_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1312_c11_6062] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_left;
     BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_return_output := BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1291_c2_f936_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1291_c6_b69f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1296_c7_c406_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1296_c11_46d4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_0719_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1303_c11_4403_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1312_c11_6062_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c11_1342_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1300_l1304_DUPLICATE_a97b_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l1300_l1304_DUPLICATE_a97b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1291_l1303_l1296_l1299_DUPLICATE_8b2f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1291_l1303_l1296_l1299_DUPLICATE_8b2f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1291_l1303_l1296_l1299_DUPLICATE_8b2f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1291_l1303_l1296_l1299_DUPLICATE_8b2f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1303_l1299_l1296_l1317_l1312_DUPLICATE_f522_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1303_l1299_l1296_l1317_l1312_DUPLICATE_f522_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1303_l1299_l1296_l1317_l1312_DUPLICATE_f522_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1303_l1299_l1296_l1317_l1312_DUPLICATE_f522_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1303_l1299_l1296_l1317_l1312_DUPLICATE_f522_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_1730_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_1730_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_1730_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_1730_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1299_l1296_l1291_l1317_l1312_DUPLICATE_9bdc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1299_l1296_l1291_l1317_l1312_DUPLICATE_9bdc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1299_l1296_l1291_l1317_l1312_DUPLICATE_9bdc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1299_l1296_l1291_l1317_l1312_DUPLICATE_9bdc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1299_l1296_l1291_l1317_l1312_DUPLICATE_9bdc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1312_l1299_DUPLICATE_00f9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1312_l1299_DUPLICATE_00f9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_29dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_29dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_29dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1291_l1296_l1312_l1299_DUPLICATE_29dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1307_c30_c1ae_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1303_c7_4f8c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l1304_c3_62bd] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_left;
     BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_return_output := BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1291_c1_6d0b] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l1315_c21_ce1e] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1315_c21_ce1e_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l1315_c31_5358_return_output);

     -- CONST_SL_8[uxn_opcodes_h_l1301_c3_eebc] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc_x <= VAR_CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc_return_output := CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1317_c7_cdaf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1312_c7_755d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1312_c7_755d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1317_c7_cdaf] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output;

     -- Submodule level 2
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_left := VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l1304_c3_62bd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1315_c21_ce1e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l1301_c3_eebc_return_output;
     VAR_printf_uxn_opcodes_h_l1292_c3_5656_uxn_opcodes_h_l1292_c3_5656_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1291_c1_6d0b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1312_c7_755d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c7_cdaf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1312_c7_755d_return_output;
     -- t16_MUX[uxn_opcodes_h_l1303_c7_4f8c] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond <= VAR_t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond;
     t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue;
     t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output := t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1305_c11_9b82] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1303_c7_4f8c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1299_c7_0cc4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;

     -- printf_uxn_opcodes_h_l1292_c3_5656[uxn_opcodes_h_l1292_c3_5656] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1292_c3_5656_uxn_opcodes_h_l1292_c3_5656_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1292_c3_5656_uxn_opcodes_h_l1292_c3_5656_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1312_c7_755d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1312_c7_755d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1312_c7_755d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1303_c7_4f8c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;

     -- Submodule level 3
     VAR_tmp16_uxn_opcodes_h_l1305_c3_7ebe := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1305_c11_9b82_return_output, 16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1312_c7_755d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1312_c7_755d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1312_c7_755d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue := VAR_tmp16_uxn_opcodes_h_l1305_c3_7ebe;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1296_c7_c406] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1303_c7_4f8c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;

     -- t16_MUX[uxn_opcodes_h_l1299_c7_0cc4] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond <= VAR_t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond;
     t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue;
     t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output := t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1299_c7_0cc4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1303_c7_4f8c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1299_c7_0cc4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1303_c7_4f8c] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond;
     tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output := tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l1310_c21_2ef9] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1310_c21_2ef9_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_tmp16_uxn_opcodes_h_l1305_c3_7ebe);

     -- Submodule level 4
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l1310_c21_2ef9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1303_c7_4f8c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1291_c2_f936] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1296_c7_c406] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1296_c7_c406] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1299_c7_0cc4] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond;
     tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output := tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;

     -- t16_MUX[uxn_opcodes_h_l1296_c7_c406] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1296_c7_c406_cond <= VAR_t16_MUX_uxn_opcodes_h_l1296_c7_c406_cond;
     t16_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue;
     t16_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output := t16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1299_c7_0cc4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1299_c7_0cc4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1303_c7_4f8c_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;
     -- t16_MUX[uxn_opcodes_h_l1291_c2_f936] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1291_c2_f936_cond <= VAR_t16_MUX_uxn_opcodes_h_l1291_c2_f936_cond;
     t16_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue;
     t16_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output := t16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1291_c2_f936] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1296_c7_c406] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_cond;
     tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output := tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1296_c7_c406] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1299_c7_0cc4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1296_c7_c406] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1291_c2_f936] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1299_c7_0cc4_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1291_c2_f936] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1296_c7_c406] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_return_output := result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1291_c2_f936] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1291_c2_f936] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_cond;
     tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output := tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output;

     -- Submodule level 7
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1296_c7_c406_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l1291_c2_f936_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1291_c2_f936] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_return_output := result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1322_l1287_DUPLICATE_4025 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1322_l1287_DUPLICATE_4025_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8c29(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1291_c2_f936_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1291_c2_f936_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1291_c2_f936_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1291_c2_f936_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1291_c2_f936_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1322_l1287_DUPLICATE_4025_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1322_l1287_DUPLICATE_4025_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
