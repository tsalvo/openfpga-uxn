-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity inc_0CLK_17cc5023 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc_0CLK_17cc5023;
architecture arch of inc_0CLK_17cc5023 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1437_c6_36aa]
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1437_c2_b835]
signal t8_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1437_c2_b835]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1437_c2_b835]
signal result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1437_c2_b835]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1437_c2_b835]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1437_c2_b835]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1437_c2_b835]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1442_c11_7a38]
signal BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1442_c7_ae2d]
signal t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1442_c7_ae2d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1442_c7_ae2d]
signal result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1442_c7_ae2d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1442_c7_ae2d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1442_c7_ae2d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1442_c7_ae2d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1445_c11_adde]
signal BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1445_c7_f447]
signal t8_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1445_c7_f447]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1445_c7_f447]
signal result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1445_c7_f447]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1445_c7_f447]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1445_c7_f447]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1445_c7_f447]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1448_c32_3b43]
signal BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1448_c32_2ece]
signal BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1448_c32_dc89]
signal MUX_uxn_opcodes_h_l1448_c32_dc89_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1448_c32_dc89_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1448_c32_dc89_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1448_c32_dc89_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1450_c11_7a3d]
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1450_c7_15b6]
signal result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1450_c7_15b6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1450_c7_15b6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1450_c7_15b6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1450_c7_15b6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1454_c24_788b]
signal BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1456_c11_f398]
signal BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1456_c7_f179]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1456_c7_f179]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_value := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_opc_done := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_left,
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_right,
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_return_output);

-- t8_MUX_uxn_opcodes_h_l1437_c2_b835
t8_MUX_uxn_opcodes_h_l1437_c2_b835 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1437_c2_b835_cond,
t8_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue,
t8_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse,
t8_MUX_uxn_opcodes_h_l1437_c2_b835_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835
result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_cond,
result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835
result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38
BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_left,
BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_right,
BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_return_output);

-- t8_MUX_uxn_opcodes_h_l1442_c7_ae2d
t8_MUX_uxn_opcodes_h_l1442_c7_ae2d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond,
t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue,
t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse,
t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d
result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond,
result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d
result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d
result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d
result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde
BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_left,
BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_right,
BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_return_output);

-- t8_MUX_uxn_opcodes_h_l1445_c7_f447
t8_MUX_uxn_opcodes_h_l1445_c7_f447 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1445_c7_f447_cond,
t8_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue,
t8_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse,
t8_MUX_uxn_opcodes_h_l1445_c7_f447_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447
result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447
result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_cond,
result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447
result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447
result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447
result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43
BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_left,
BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_right,
BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece
BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_left,
BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_right,
BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_return_output);

-- MUX_uxn_opcodes_h_l1448_c32_dc89
MUX_uxn_opcodes_h_l1448_c32_dc89 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1448_c32_dc89_cond,
MUX_uxn_opcodes_h_l1448_c32_dc89_iftrue,
MUX_uxn_opcodes_h_l1448_c32_dc89_iffalse,
MUX_uxn_opcodes_h_l1448_c32_dc89_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_left,
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_right,
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6
result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_cond,
result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6
result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b
BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_left,
BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_right,
BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398
BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_left,
BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_right,
BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179
result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179
result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_return_output,
 t8_MUX_uxn_opcodes_h_l1437_c2_b835_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_return_output,
 t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_return_output,
 t8_MUX_uxn_opcodes_h_l1445_c7_f447_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_return_output,
 MUX_uxn_opcodes_h_l1448_c32_dc89_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1439_c3_4fa9 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1443_c3_062d : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1448_c32_dc89_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1448_c32_dc89_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1448_c32_dc89_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1448_c32_dc89_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_uxn_opcodes_h_l1454_c3_0e9d : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1453_c3_ba9c : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_return_output : unsigned(8 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1442_l1445_l1437_DUPLICATE_23a6_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1442_l1445_l1437_l1450_DUPLICATE_ed78_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1442_l1437_l1450_DUPLICATE_41cc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_8525_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1450_DUPLICATE_ceae_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1445_l1450_DUPLICATE_8004_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l1461_l1433_DUPLICATE_4a51_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1443_c3_062d := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1443_c3_062d;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_right := to_unsigned(3, 2);
     VAR_MUX_uxn_opcodes_h_l1448_c32_dc89_iffalse := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_right := to_unsigned(1, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_right := to_unsigned(128, 8);
     VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_right := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1448_c32_dc89_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1453_c3_ba9c := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1453_c3_ba9c;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1439_c3_4fa9 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1439_c3_4fa9;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_right := to_unsigned(0, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse := t8;
     -- BIN_OP_PLUS[uxn_opcodes_h_l1454_c24_788b] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1442_l1445_l1437_l1450_DUPLICATE_ed78 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1442_l1445_l1437_l1450_DUPLICATE_ed78_return_output := result.stack_value;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1442_l1445_l1437_DUPLICATE_23a6 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1442_l1445_l1437_DUPLICATE_23a6_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1450_c11_7a3d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1445_c11_adde] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_left;
     BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_return_output := BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1456_c11_f398] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_left;
     BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_return_output := BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1445_l1450_DUPLICATE_8004 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1445_l1450_DUPLICATE_8004_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1437_c6_36aa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_left;
     BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_return_output := BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_8525 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_8525_return_output := result.is_stack_write;

     -- BIN_OP_AND[uxn_opcodes_h_l1448_c32_3b43] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_left;
     BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_return_output := BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1442_l1437_l1450_DUPLICATE_41cc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1442_l1437_l1450_DUPLICATE_41cc_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1450_DUPLICATE_ceae LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1450_DUPLICATE_ceae_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1442_c11_7a38] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_left;
     BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_return_output := BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_3b43_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_b835_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_36aa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_7a38_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1445_c7_f447_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_adde_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_7a3d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_f398_return_output;
     VAR_result_stack_value_uxn_opcodes_h_l1454_c3_0e9d := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_788b_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1442_l1445_l1437_DUPLICATE_23a6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1442_l1445_l1437_DUPLICATE_23a6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1442_l1445_l1437_DUPLICATE_23a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1450_DUPLICATE_ceae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1450_DUPLICATE_ceae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1450_DUPLICATE_ceae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1450_DUPLICATE_ceae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1442_l1437_l1450_DUPLICATE_41cc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1442_l1437_l1450_DUPLICATE_41cc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1442_l1437_l1450_DUPLICATE_41cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_8525_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_8525_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_8525_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_8525_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1445_l1450_DUPLICATE_8004_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1445_l1450_DUPLICATE_8004_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1442_l1445_l1437_l1450_DUPLICATE_ed78_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1442_l1445_l1437_l1450_DUPLICATE_ed78_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1442_l1445_l1437_l1450_DUPLICATE_ed78_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1442_l1445_l1437_l1450_DUPLICATE_ed78_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue := VAR_result_stack_value_uxn_opcodes_h_l1454_c3_0e9d;
     -- result_stack_value_MUX[uxn_opcodes_h_l1450_c7_15b6] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output := result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1450_c7_15b6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1456_c7_f179] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1448_c32_2ece] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_left;
     BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_return_output := BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_return_output;

     -- t8_MUX[uxn_opcodes_h_l1445_c7_f447] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1445_c7_f447_cond <= VAR_t8_MUX_uxn_opcodes_h_l1445_c7_f447_cond;
     t8_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue;
     t8_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1445_c7_f447_return_output := t8_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1456_c7_f179] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1450_c7_15b6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1448_c32_dc89_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_2ece_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_f179_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_f179_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1445_c7_f447] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1445_c7_f447] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_return_output := result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;

     -- MUX[uxn_opcodes_h_l1448_c32_dc89] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1448_c32_dc89_cond <= VAR_MUX_uxn_opcodes_h_l1448_c32_dc89_cond;
     MUX_uxn_opcodes_h_l1448_c32_dc89_iftrue <= VAR_MUX_uxn_opcodes_h_l1448_c32_dc89_iftrue;
     MUX_uxn_opcodes_h_l1448_c32_dc89_iffalse <= VAR_MUX_uxn_opcodes_h_l1448_c32_dc89_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1448_c32_dc89_return_output := MUX_uxn_opcodes_h_l1448_c32_dc89_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1450_c7_15b6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output;

     -- t8_MUX[uxn_opcodes_h_l1442_c7_ae2d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond <= VAR_t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond;
     t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue;
     t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output := t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1445_c7_f447] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1450_c7_15b6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue := VAR_MUX_uxn_opcodes_h_l1448_c32_dc89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_15b6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1445_c7_f447] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1442_c7_ae2d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1442_c7_ae2d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1445_c7_f447] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1442_c7_ae2d] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output := result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;

     -- t8_MUX[uxn_opcodes_h_l1437_c2_b835] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1437_c2_b835_cond <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_b835_cond;
     t8_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue;
     t8_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_b835_return_output := t8_MUX_uxn_opcodes_h_l1437_c2_b835_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1445_c7_f447] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_f447_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1437_c2_b835_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1437_c2_b835] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1437_c2_b835] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_return_output := result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1442_c7_ae2d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1442_c7_ae2d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1442_c7_ae2d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1437_c2_b835] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_ae2d_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1437_c2_b835] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1437_c2_b835] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1437_c2_b835] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l1461_l1433_DUPLICATE_4a51 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l1461_l1433_DUPLICATE_4a51_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_b835_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_b835_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_b835_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_b835_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_b835_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l1461_l1433_DUPLICATE_4a51_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l1461_l1433_DUPLICATE_4a51_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
