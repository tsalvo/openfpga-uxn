-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 57
entity opc_deo_phased_0CLK_1b2abcad is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_deo_phased_0CLK_1b2abcad;
architecture arch of opc_deo_phased_0CLK_1b2abcad is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l912_c6_4042]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l912_c1_30f9]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l916_c7_b979]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l912_c2_e3a5]
signal t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l912_c2_e3a5]
signal n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l912_c2_e3a5]
signal result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output : unsigned(0 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l913_c12_18e5]
signal set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_return_output : unsigned(0 downto 0);

-- t_register[uxn_opcodes_phased_h_l914_c8_0522]
signal t_register_uxn_opcodes_phased_h_l914_c8_0522_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l914_c8_0522_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l914_c8_0522_stack_ptr : unsigned(7 downto 0);
signal t_register_uxn_opcodes_phased_h_l914_c8_0522_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l916_c11_1eb7]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l916_c1_4b31]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l919_c7_ae4b]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l916_c7_b979]
signal t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l916_c7_b979]
signal n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l916_c7_b979]
signal result_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l917_c8_8204]
signal n_register_uxn_opcodes_phased_h_l917_c8_8204_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l917_c8_8204_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l917_c8_8204_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l917_c8_8204_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l919_c11_aba0]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l919_c1_31fb]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l922_c7_6c25]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l919_c7_ae4b]
signal n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l919_c7_ae4b]
signal result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l920_c8_3ec6]
signal n_register_uxn_opcodes_phased_h_l920_c8_3ec6_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l920_c8_3ec6_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l920_c8_3ec6_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l920_c8_3ec6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l922_c11_0698]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l922_c1_f4b6]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l925_c7_5c40]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l922_c7_6c25]
signal result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output : unsigned(0 downto 0);

-- set[uxn_opcodes_phased_h_l923_c3_c35a]
signal set_uxn_opcodes_phased_h_l923_c3_c35a_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l923_c3_c35a_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l923_c3_c35a_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l923_c3_c35a_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l923_c3_c35a_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l923_c3_c35a_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l923_c3_c35a_add : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l925_c11_99cc]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l925_c1_ec03]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l928_c7_264c]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l925_c7_5c40]
signal result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output : unsigned(0 downto 0);

-- deo_phased[uxn_opcodes_phased_h_l926_c12_cd4c]
signal deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_CLOCK_ENABLE : unsigned(0 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_phase : unsigned(3 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_device_address : unsigned(7 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_value : unsigned(7 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l928_c11_0815]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l928_c1_4785]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l931_c7_fe48]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l928_c7_264c]
signal result_MUX_uxn_opcodes_phased_h_l928_c7_264c_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l928_c7_264c_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l928_c7_264c_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output : unsigned(0 downto 0);

-- deo_phased[uxn_opcodes_phased_h_l929_c12_5530]
signal deo_phased_uxn_opcodes_phased_h_l929_c12_5530_CLOCK_ENABLE : unsigned(0 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l929_c12_5530_phase : unsigned(3 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l929_c12_5530_device_address : unsigned(7 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l929_c12_5530_value : unsigned(7 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l929_c12_5530_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l931_c11_a9a6]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l931_c1_5152]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l934_c7_8d56]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l931_c7_fe48]
signal result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output : unsigned(0 downto 0);

-- deo_phased[uxn_opcodes_phased_h_l932_c12_3387]
signal deo_phased_uxn_opcodes_phased_h_l932_c12_3387_CLOCK_ENABLE : unsigned(0 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l932_c12_3387_phase : unsigned(3 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l932_c12_3387_device_address : unsigned(7 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l932_c12_3387_value : unsigned(7 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l932_c12_3387_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l934_c11_b47f]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l934_c1_0c58]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l937_c7_cabd]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l934_c7_8d56]
signal result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output : unsigned(0 downto 0);

-- deo_phased[uxn_opcodes_phased_h_l935_c12_d0a8]
signal deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_CLOCK_ENABLE : unsigned(0 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_phase : unsigned(3 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_device_address : unsigned(7 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_value : unsigned(7 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l937_c11_20b8]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_right : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l937_c1_a291]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l940_c7_e3a6]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l937_c7_cabd]
signal result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output : unsigned(0 downto 0);

-- deo_phased[uxn_opcodes_phased_h_l938_c12_50e3]
signal deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_CLOCK_ENABLE : unsigned(0 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_phase : unsigned(3 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_device_address : unsigned(7 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_value : unsigned(7 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l940_c11_9b3b]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_right : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l940_c1_5397]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l940_c7_e3a6]
signal result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output : unsigned(0 downto 0);

-- deo_phased[uxn_opcodes_phased_h_l941_c12_5abf]
signal deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_CLOCK_ENABLE : unsigned(0 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_phase : unsigned(3 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_device_address : unsigned(7 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_value : unsigned(7 downto 0);
signal deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l943_c11_3fb0]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_right : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l943_c7_e347]
signal result_MUX_uxn_opcodes_phased_h_l943_c7_e347_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l943_c7_e347_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l943_c7_e347_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l943_c7_e347_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042
BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5
t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond,
t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue,
t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse,
t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5
n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond,
n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue,
n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse,
n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output);

-- result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5
result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond,
result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue,
result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse,
result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5
set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5 : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_sp,
set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_k,
set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_mul,
set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_add,
set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_return_output);

-- t_register_uxn_opcodes_phased_h_l914_c8_0522
t_register_uxn_opcodes_phased_h_l914_c8_0522 : entity work.t_register_0CLK_621d5f60 port map (
clk,
t_register_uxn_opcodes_phased_h_l914_c8_0522_CLOCK_ENABLE,
t_register_uxn_opcodes_phased_h_l914_c8_0522_stack_index,
t_register_uxn_opcodes_phased_h_l914_c8_0522_stack_ptr,
t_register_uxn_opcodes_phased_h_l914_c8_0522_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7
BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l916_c7_b979
t8_MUX_uxn_opcodes_phased_h_l916_c7_b979 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond,
t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue,
t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse,
t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l916_c7_b979
n8_MUX_uxn_opcodes_phased_h_l916_c7_b979 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond,
n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue,
n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse,
n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output);

-- result_MUX_uxn_opcodes_phased_h_l916_c7_b979
result_MUX_uxn_opcodes_phased_h_l916_c7_b979 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond,
result_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue,
result_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse,
result_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output);

-- n_register_uxn_opcodes_phased_h_l917_c8_8204
n_register_uxn_opcodes_phased_h_l917_c8_8204 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l917_c8_8204_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l917_c8_8204_stack_index,
n_register_uxn_opcodes_phased_h_l917_c8_8204_stack_ptr,
n_register_uxn_opcodes_phased_h_l917_c8_8204_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0
BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b
n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond,
n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue,
n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse,
n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output);

-- result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b
result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond,
result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue,
result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse,
result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output);

-- n_register_uxn_opcodes_phased_h_l920_c8_3ec6
n_register_uxn_opcodes_phased_h_l920_c8_3ec6 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l920_c8_3ec6_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l920_c8_3ec6_stack_index,
n_register_uxn_opcodes_phased_h_l920_c8_3ec6_stack_ptr,
n_register_uxn_opcodes_phased_h_l920_c8_3ec6_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698
BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output);

-- result_MUX_uxn_opcodes_phased_h_l922_c7_6c25
result_MUX_uxn_opcodes_phased_h_l922_c7_6c25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_cond,
result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iftrue,
result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iffalse,
result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output);

-- set_uxn_opcodes_phased_h_l923_c3_c35a
set_uxn_opcodes_phased_h_l923_c3_c35a : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l923_c3_c35a_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l923_c3_c35a_sp,
set_uxn_opcodes_phased_h_l923_c3_c35a_stack_index,
set_uxn_opcodes_phased_h_l923_c3_c35a_ins,
set_uxn_opcodes_phased_h_l923_c3_c35a_k,
set_uxn_opcodes_phased_h_l923_c3_c35a_mul,
set_uxn_opcodes_phased_h_l923_c3_c35a_add);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc
BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output);

-- result_MUX_uxn_opcodes_phased_h_l925_c7_5c40
result_MUX_uxn_opcodes_phased_h_l925_c7_5c40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_cond,
result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iftrue,
result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iffalse,
result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output);

-- deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c
deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c : entity work.deo_phased_0CLK_0ef75794 port map (
clk,
deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_CLOCK_ENABLE,
deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_phase,
deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_device_address,
deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_value,
deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815
BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output);

-- result_MUX_uxn_opcodes_phased_h_l928_c7_264c
result_MUX_uxn_opcodes_phased_h_l928_c7_264c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l928_c7_264c_cond,
result_MUX_uxn_opcodes_phased_h_l928_c7_264c_iftrue,
result_MUX_uxn_opcodes_phased_h_l928_c7_264c_iffalse,
result_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output);

-- deo_phased_uxn_opcodes_phased_h_l929_c12_5530
deo_phased_uxn_opcodes_phased_h_l929_c12_5530 : entity work.deo_phased_0CLK_0ef75794 port map (
clk,
deo_phased_uxn_opcodes_phased_h_l929_c12_5530_CLOCK_ENABLE,
deo_phased_uxn_opcodes_phased_h_l929_c12_5530_phase,
deo_phased_uxn_opcodes_phased_h_l929_c12_5530_device_address,
deo_phased_uxn_opcodes_phased_h_l929_c12_5530_value,
deo_phased_uxn_opcodes_phased_h_l929_c12_5530_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6
BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output);

-- result_MUX_uxn_opcodes_phased_h_l931_c7_fe48
result_MUX_uxn_opcodes_phased_h_l931_c7_fe48 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_cond,
result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iftrue,
result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iffalse,
result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output);

-- deo_phased_uxn_opcodes_phased_h_l932_c12_3387
deo_phased_uxn_opcodes_phased_h_l932_c12_3387 : entity work.deo_phased_0CLK_0ef75794 port map (
clk,
deo_phased_uxn_opcodes_phased_h_l932_c12_3387_CLOCK_ENABLE,
deo_phased_uxn_opcodes_phased_h_l932_c12_3387_phase,
deo_phased_uxn_opcodes_phased_h_l932_c12_3387_device_address,
deo_phased_uxn_opcodes_phased_h_l932_c12_3387_value,
deo_phased_uxn_opcodes_phased_h_l932_c12_3387_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f
BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output);

-- result_MUX_uxn_opcodes_phased_h_l934_c7_8d56
result_MUX_uxn_opcodes_phased_h_l934_c7_8d56 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_cond,
result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iftrue,
result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iffalse,
result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output);

-- deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8
deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8 : entity work.deo_phased_0CLK_0ef75794 port map (
clk,
deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_CLOCK_ENABLE,
deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_phase,
deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_device_address,
deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_value,
deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8
BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output);

-- result_MUX_uxn_opcodes_phased_h_l937_c7_cabd
result_MUX_uxn_opcodes_phased_h_l937_c7_cabd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_cond,
result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iftrue,
result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iffalse,
result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output);

-- deo_phased_uxn_opcodes_phased_h_l938_c12_50e3
deo_phased_uxn_opcodes_phased_h_l938_c12_50e3 : entity work.deo_phased_0CLK_0ef75794 port map (
clk,
deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_CLOCK_ENABLE,
deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_phase,
deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_device_address,
deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_value,
deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b
BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_return_output);

-- result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6
result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_cond,
result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iftrue,
result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iffalse,
result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output);

-- deo_phased_uxn_opcodes_phased_h_l941_c12_5abf
deo_phased_uxn_opcodes_phased_h_l941_c12_5abf : entity work.deo_phased_0CLK_0ef75794 port map (
clk,
deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_CLOCK_ENABLE,
deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_phase,
deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_device_address,
deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_value,
deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0
BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_return_output);

-- result_MUX_uxn_opcodes_phased_h_l943_c7_e347
result_MUX_uxn_opcodes_phased_h_l943_c7_e347 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l943_c7_e347_cond,
result_MUX_uxn_opcodes_phased_h_l943_c7_e347_iftrue,
result_MUX_uxn_opcodes_phased_h_l943_c7_e347_iffalse,
result_MUX_uxn_opcodes_phased_h_l943_c7_e347_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 n8,
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output,
 t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output,
 n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output,
 result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output,
 set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_return_output,
 t_register_uxn_opcodes_phased_h_l914_c8_0522_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output,
 t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output,
 n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output,
 result_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output,
 n_register_uxn_opcodes_phased_h_l917_c8_8204_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output,
 n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output,
 result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output,
 n_register_uxn_opcodes_phased_h_l920_c8_3ec6_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output,
 result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output,
 result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output,
 deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output,
 result_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output,
 deo_phased_uxn_opcodes_phased_h_l929_c12_5530_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output,
 result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output,
 deo_phased_uxn_opcodes_phased_h_l932_c12_3387_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output,
 result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output,
 deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output,
 result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output,
 deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_return_output,
 result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output,
 deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_return_output,
 result_MUX_uxn_opcodes_phased_h_l943_c7_e347_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_return_output : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l914_c8_0522_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l914_c8_0522_stack_ptr : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l914_c8_0522_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l914_c8_0522_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l917_c8_8204_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l917_c8_8204_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l917_c8_8204_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l917_c8_8204_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l920_c8_3ec6_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l920_c8_3ec6_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l920_c8_3ec6_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l920_c8_3ec6_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_cond : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_cond : unsigned(0 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_phase : unsigned(3 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_device_address : unsigned(7 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_value : unsigned(7 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l928_c7_264c_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l928_c7_264c_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l928_c7_264c_cond : unsigned(0 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_phase : unsigned(3 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_device_address : unsigned(7 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_value : unsigned(7 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_cond : unsigned(0 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_phase : unsigned(3 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_device_address : unsigned(7 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_value : unsigned(7 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_cond : unsigned(0 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_phase : unsigned(3 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_device_address : unsigned(7 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_value : unsigned(7 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_cond : unsigned(0 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_phase : unsigned(3 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_device_address : unsigned(7 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_value : unsigned(7 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l943_c7_e347_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_cond : unsigned(0 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_phase : unsigned(3 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_device_address : unsigned(7 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_value : unsigned(7 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l943_c7_e347_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l943_c7_e347_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l943_c7_e347_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_n8 := n8;
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_right := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_right := to_unsigned(9, 4);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_right := to_unsigned(3, 2);
     VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_phase := resize(to_unsigned(5, 3), 4);
     VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_add := resize(to_signed(-2, 3), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue := to_unsigned(0, 1);
     VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_phase := resize(to_unsigned(0, 1), 4);
     VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_add := resize(to_signed(-2, 3), 8);
     VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_phase := resize(to_unsigned(2, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_right := to_unsigned(8, 4);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_right := to_unsigned(7, 3);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_iffalse := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_right := to_unsigned(6, 3);
     VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_phase := resize(to_unsigned(3, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iftrue := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_iffalse := to_unsigned(0, 1);
     VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_mul := resize(to_unsigned(2, 2), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_iffalse := to_unsigned(0, 1);
     VAR_result_MUX_uxn_opcodes_phased_h_l943_c7_e347_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_right := to_unsigned(10, 4);
     VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_phase := resize(to_unsigned(4, 3), 4);
     VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_phase := resize(to_unsigned(1, 1), 4);
     VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_mul := resize(to_unsigned(2, 2), 8);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_iffalse := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_k := VAR_k;
     VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_value := n8;
     VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_value := n8;
     VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_value := n8;
     VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_value := n8;
     VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_value := n8;
     VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_value := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_left := VAR_phase;
     VAR_result_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l943_c7_e347_iffalse := result;
     VAR_n_register_uxn_opcodes_phased_h_l917_c8_8204_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l920_c8_3ec6_stack_ptr := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_sp := VAR_sp;
     VAR_t_register_uxn_opcodes_phased_h_l914_c8_0522_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l917_c8_8204_stack_index := VAR_stack_index;
     VAR_n_register_uxn_opcodes_phased_h_l920_c8_3ec6_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_phased_h_l914_c8_0522_stack_index := VAR_stack_index;
     VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_device_address := t8;
     VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_device_address := t8;
     VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_device_address := t8;
     VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_device_address := t8;
     VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_device_address := t8;
     VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_device_address := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_phased_h_l931_c11_a9a6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l940_c11_9b3b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l916_c11_1eb7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l919_c11_aba0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l937_c11_20b8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l934_c11_b47f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l928_c11_0815] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l943_c11_3fb0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l925_c11_99cc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l912_c6_4042] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l922_c11_0698] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l912_c6_4042_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l916_c11_1eb7_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l919_c11_aba0_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l922_c11_0698_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l925_c11_99cc_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l928_c7_264c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l928_c11_0815_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l931_c11_a9a6_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l934_c11_b47f_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l937_c11_20b8_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l940_c11_9b3b_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l943_c7_e347_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l943_c11_3fb0_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l916_c7_b979] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l912_c1_30f9] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l943_c7_e347] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l943_c7_e347_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l943_c7_e347_cond;
     result_MUX_uxn_opcodes_phased_h_l943_c7_e347_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l943_c7_e347_iftrue;
     result_MUX_uxn_opcodes_phased_h_l943_c7_e347_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l943_c7_e347_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l943_c7_e347_return_output := result_MUX_uxn_opcodes_phased_h_l943_c7_e347_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_return_output;
     VAR_t_register_uxn_opcodes_phased_h_l914_c8_0522_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l912_c1_30f9_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l943_c7_e347_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l919_c7_ae4b] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l916_c1_4b31] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_return_output;

     -- t_register[uxn_opcodes_phased_h_l914_c8_0522] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_phased_h_l914_c8_0522_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_phased_h_l914_c8_0522_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_phased_h_l914_c8_0522_stack_index <= VAR_t_register_uxn_opcodes_phased_h_l914_c8_0522_stack_index;
     t_register_uxn_opcodes_phased_h_l914_c8_0522_stack_ptr <= VAR_t_register_uxn_opcodes_phased_h_l914_c8_0522_stack_ptr;
     -- Outputs
     VAR_t_register_uxn_opcodes_phased_h_l914_c8_0522_return_output := t_register_uxn_opcodes_phased_h_l914_c8_0522_return_output;

     -- set_will_fail[uxn_opcodes_phased_h_l913_c12_18e5] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_sp;
     set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_k;
     set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_mul;
     set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_return_output := set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l917_c8_8204_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l916_c1_4b31_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l913_c12_18e5_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue := VAR_t_register_uxn_opcodes_phased_h_l914_c8_0522_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l922_c7_6c25] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output;

     -- n_register[uxn_opcodes_phased_h_l917_c8_8204] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l917_c8_8204_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l917_c8_8204_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l917_c8_8204_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l917_c8_8204_stack_index;
     n_register_uxn_opcodes_phased_h_l917_c8_8204_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l917_c8_8204_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l917_c8_8204_return_output := n_register_uxn_opcodes_phased_h_l917_c8_8204_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l919_c1_31fb] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l920_c8_3ec6_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l919_c1_31fb_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue := VAR_n_register_uxn_opcodes_phased_h_l917_c8_8204_return_output;
     -- n_register[uxn_opcodes_phased_h_l920_c8_3ec6] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l920_c8_3ec6_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l920_c8_3ec6_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l920_c8_3ec6_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l920_c8_3ec6_stack_index;
     n_register_uxn_opcodes_phased_h_l920_c8_3ec6_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l920_c8_3ec6_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l920_c8_3ec6_return_output := n_register_uxn_opcodes_phased_h_l920_c8_3ec6_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l922_c1_f4b6] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l916_c7_b979] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond;
     t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output := t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l925_c7_5c40] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output;

     -- Submodule level 5
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output;
     VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l922_c1_f4b6_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue := VAR_n_register_uxn_opcodes_phased_h_l920_c8_3ec6_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output;
     -- t8_MUX[uxn_opcodes_phased_h_l912_c2_e3a5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond;
     t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output := t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l928_c7_264c] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l925_c1_ec03] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_return_output;

     -- n8_MUX[uxn_opcodes_phased_h_l919_c7_ae4b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond;
     n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output := n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output;

     -- set[uxn_opcodes_phased_h_l923_c3_c35a] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l923_c3_c35a_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l923_c3_c35a_sp <= VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_sp;
     set_uxn_opcodes_phased_h_l923_c3_c35a_stack_index <= VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_stack_index;
     set_uxn_opcodes_phased_h_l923_c3_c35a_ins <= VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_ins;
     set_uxn_opcodes_phased_h_l923_c3_c35a_k <= VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_k;
     set_uxn_opcodes_phased_h_l923_c3_c35a_mul <= VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_mul;
     set_uxn_opcodes_phased_h_l923_c3_c35a_add <= VAR_set_uxn_opcodes_phased_h_l923_c3_c35a_add;
     -- Outputs

     -- Submodule level 6
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output;
     VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l925_c1_ec03_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l928_c1_4785] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_return_output;

     -- n8_MUX[uxn_opcodes_phased_h_l916_c7_b979] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond;
     n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output := n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l931_c7_fe48] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output;

     -- deo_phased[uxn_opcodes_phased_h_l926_c12_cd4c] LATENCY=0
     -- Clock enable
     deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_CLOCK_ENABLE <= VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_CLOCK_ENABLE;
     -- Inputs
     deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_phase <= VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_phase;
     deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_device_address <= VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_device_address;
     deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_value <= VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_value;
     -- Outputs
     VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_return_output := deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_return_output;

     -- Submodule level 7
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output;
     VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l928_c1_4785_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iftrue := VAR_deo_phased_uxn_opcodes_phased_h_l926_c12_cd4c_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l912_c2_e3a5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond;
     n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output := n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output;

     -- deo_phased[uxn_opcodes_phased_h_l929_c12_5530] LATENCY=0
     -- Clock enable
     deo_phased_uxn_opcodes_phased_h_l929_c12_5530_CLOCK_ENABLE <= VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_CLOCK_ENABLE;
     -- Inputs
     deo_phased_uxn_opcodes_phased_h_l929_c12_5530_phase <= VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_phase;
     deo_phased_uxn_opcodes_phased_h_l929_c12_5530_device_address <= VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_device_address;
     deo_phased_uxn_opcodes_phased_h_l929_c12_5530_value <= VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_value;
     -- Outputs
     VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_return_output := deo_phased_uxn_opcodes_phased_h_l929_c12_5530_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l931_c1_5152] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l934_c7_8d56] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output;

     -- Submodule level 8
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output;
     VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l931_c1_5152_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l928_c7_264c_iftrue := VAR_deo_phased_uxn_opcodes_phased_h_l929_c12_5530_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l937_c7_cabd] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l934_c1_0c58] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_return_output;

     -- deo_phased[uxn_opcodes_phased_h_l932_c12_3387] LATENCY=0
     -- Clock enable
     deo_phased_uxn_opcodes_phased_h_l932_c12_3387_CLOCK_ENABLE <= VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_CLOCK_ENABLE;
     -- Inputs
     deo_phased_uxn_opcodes_phased_h_l932_c12_3387_phase <= VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_phase;
     deo_phased_uxn_opcodes_phased_h_l932_c12_3387_device_address <= VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_device_address;
     deo_phased_uxn_opcodes_phased_h_l932_c12_3387_value <= VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_value;
     -- Outputs
     VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_return_output := deo_phased_uxn_opcodes_phased_h_l932_c12_3387_return_output;

     -- Submodule level 9
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output;
     VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l934_c1_0c58_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iftrue := VAR_deo_phased_uxn_opcodes_phased_h_l932_c12_3387_return_output;
     -- deo_phased[uxn_opcodes_phased_h_l935_c12_d0a8] LATENCY=0
     -- Clock enable
     deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_CLOCK_ENABLE <= VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_CLOCK_ENABLE;
     -- Inputs
     deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_phase <= VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_phase;
     deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_device_address <= VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_device_address;
     deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_value <= VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_value;
     -- Outputs
     VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_return_output := deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l937_c1_a291] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l940_c7_e3a6] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output;

     -- Submodule level 10
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output;
     VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l937_c1_a291_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iftrue := VAR_deo_phased_uxn_opcodes_phased_h_l935_c12_d0a8_return_output;
     -- deo_phased[uxn_opcodes_phased_h_l938_c12_50e3] LATENCY=0
     -- Clock enable
     deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_CLOCK_ENABLE <= VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_CLOCK_ENABLE;
     -- Inputs
     deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_phase <= VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_phase;
     deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_device_address <= VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_device_address;
     deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_value <= VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_value;
     -- Outputs
     VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_return_output := deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l940_c1_5397] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_return_output;

     -- Submodule level 11
     VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l940_c1_5397_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iftrue := VAR_deo_phased_uxn_opcodes_phased_h_l938_c12_50e3_return_output;
     -- deo_phased[uxn_opcodes_phased_h_l941_c12_5abf] LATENCY=0
     -- Clock enable
     deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_CLOCK_ENABLE <= VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_CLOCK_ENABLE;
     -- Inputs
     deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_phase <= VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_phase;
     deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_device_address <= VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_device_address;
     deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_value <= VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_value;
     -- Outputs
     VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_return_output := deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_return_output;

     -- Submodule level 12
     VAR_result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iftrue := VAR_deo_phased_uxn_opcodes_phased_h_l941_c12_5abf_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l940_c7_e3a6] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_cond;
     result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iftrue;
     result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output := result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output;

     -- Submodule level 13
     VAR_result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l940_c7_e3a6_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l937_c7_cabd] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_cond;
     result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iftrue;
     result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output := result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output;

     -- Submodule level 14
     VAR_result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l937_c7_cabd_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l934_c7_8d56] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_cond;
     result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iftrue;
     result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output := result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output;

     -- Submodule level 15
     VAR_result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l934_c7_8d56_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l931_c7_fe48] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_cond;
     result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iftrue;
     result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output := result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output;

     -- Submodule level 16
     VAR_result_MUX_uxn_opcodes_phased_h_l928_c7_264c_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l931_c7_fe48_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l928_c7_264c] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l928_c7_264c_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l928_c7_264c_cond;
     result_MUX_uxn_opcodes_phased_h_l928_c7_264c_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l928_c7_264c_iftrue;
     result_MUX_uxn_opcodes_phased_h_l928_c7_264c_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l928_c7_264c_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output := result_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output;

     -- Submodule level 17
     VAR_result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l928_c7_264c_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l925_c7_5c40] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_cond;
     result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iftrue;
     result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output := result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output;

     -- Submodule level 18
     VAR_result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l925_c7_5c40_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l922_c7_6c25] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_cond;
     result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iftrue;
     result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output := result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output;

     -- Submodule level 19
     VAR_result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l922_c7_6c25_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l919_c7_ae4b] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_cond;
     result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iftrue;
     result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output := result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output;

     -- Submodule level 20
     VAR_result_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l919_c7_ae4b_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l916_c7_b979] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l916_c7_b979_cond;
     result_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l916_c7_b979_iftrue;
     result_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l916_c7_b979_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output := result_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output;

     -- Submodule level 21
     VAR_result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l916_c7_b979_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l912_c2_e3a5] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_cond;
     result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iftrue;
     result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output := result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output;

     -- Submodule level 22
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l912_c2_e3a5_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     n8 <= REG_COMB_n8;
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
