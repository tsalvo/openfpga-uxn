-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity sta2_0CLK_bce25fe8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end sta2_0CLK_bce25fe8;
architecture arch of sta2_0CLK_bce25fe8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2106_c6_ed3c]
signal BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2106_c2_563f]
signal result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2106_c2_563f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2106_c2_563f]
signal result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2106_c2_563f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2106_c2_563f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2106_c2_563f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2106_c2_563f]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2106_c2_563f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l2106_c2_563f]
signal n16_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l2106_c2_563f]
signal t16_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2114_c11_f4ef]
signal BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2114_c7_4abc]
signal result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2114_c7_4abc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2114_c7_4abc]
signal result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2114_c7_4abc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2114_c7_4abc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2114_c7_4abc]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2114_c7_4abc]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2114_c7_4abc]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l2114_c7_4abc]
signal n16_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l2114_c7_4abc]
signal t16_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2117_c11_97d2]
signal BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2117_c7_d69f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2117_c7_d69f]
signal result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2117_c7_d69f]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2117_c7_d69f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2117_c7_d69f]
signal result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2117_c7_d69f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2117_c7_d69f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l2117_c7_d69f]
signal n16_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l2117_c7_d69f]
signal t16_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2121_c30_136a]
signal sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2123_c11_18fe]
signal BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2123_c7_7514]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2123_c7_7514]
signal result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2123_c7_7514]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2123_c7_7514]
signal result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2123_c7_7514]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2123_c7_7514]
signal t16_MUX_uxn_opcodes_h_l2123_c7_7514_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2123_c7_7514_return_output : unsigned(15 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l2128_c31_d706]
signal CONST_SR_8_uxn_opcodes_h_l2128_c31_d706_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l2128_c31_d706_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2130_c11_6548]
signal BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2130_c7_333b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2130_c7_333b]
signal result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2130_c7_333b]
signal result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2130_c7_333b]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l2131_c22_9913]
signal BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2134_c11_1b33]
signal BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2134_c7_a284]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2134_c7_a284]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_sp_shift := ref_toks_6;
      base.is_stack_operation_16bit := ref_toks_7;
      base.is_ram_write := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c
BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_left,
BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_right,
BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f
result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_cond,
result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f
result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f
result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f
result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f
result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_return_output);

-- n16_MUX_uxn_opcodes_h_l2106_c2_563f
n16_MUX_uxn_opcodes_h_l2106_c2_563f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2106_c2_563f_cond,
n16_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue,
n16_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse,
n16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output);

-- t16_MUX_uxn_opcodes_h_l2106_c2_563f
t16_MUX_uxn_opcodes_h_l2106_c2_563f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2106_c2_563f_cond,
t16_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue,
t16_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse,
t16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef
BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_left,
BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_right,
BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc
result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_cond,
result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc
result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc
result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_cond,
result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc
result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc
result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc
result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output);

-- n16_MUX_uxn_opcodes_h_l2114_c7_4abc
n16_MUX_uxn_opcodes_h_l2114_c7_4abc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2114_c7_4abc_cond,
n16_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue,
n16_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse,
n16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output);

-- t16_MUX_uxn_opcodes_h_l2114_c7_4abc
t16_MUX_uxn_opcodes_h_l2114_c7_4abc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2114_c7_4abc_cond,
t16_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue,
t16_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse,
t16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2
BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_left,
BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_right,
BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f
result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f
result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_cond,
result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f
result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f
result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f
result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output);

-- n16_MUX_uxn_opcodes_h_l2117_c7_d69f
n16_MUX_uxn_opcodes_h_l2117_c7_d69f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2117_c7_d69f_cond,
n16_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue,
n16_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse,
n16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output);

-- t16_MUX_uxn_opcodes_h_l2117_c7_d69f
t16_MUX_uxn_opcodes_h_l2117_c7_d69f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2117_c7_d69f_cond,
t16_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue,
t16_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse,
t16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2121_c30_136a
sp_relative_shift_uxn_opcodes_h_l2121_c30_136a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_ins,
sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_x,
sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_y,
sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe
BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_left,
BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_right,
BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514
result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514
result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_cond,
result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514
result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514
result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_cond,
result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514
result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_return_output);

-- t16_MUX_uxn_opcodes_h_l2123_c7_7514
t16_MUX_uxn_opcodes_h_l2123_c7_7514 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2123_c7_7514_cond,
t16_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue,
t16_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse,
t16_MUX_uxn_opcodes_h_l2123_c7_7514_return_output);

-- CONST_SR_8_uxn_opcodes_h_l2128_c31_d706
CONST_SR_8_uxn_opcodes_h_l2128_c31_d706 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l2128_c31_d706_x,
CONST_SR_8_uxn_opcodes_h_l2128_c31_d706_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548
BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_left,
BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_right,
BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b
result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b
result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b
result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_cond,
result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b
result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913
BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913 : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_left,
BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_right,
BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33
BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_left,
BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_right,
BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284
result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284
result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
 n16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
 t16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output,
 n16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output,
 t16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output,
 n16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output,
 t16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output,
 sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_return_output,
 t16_MUX_uxn_opcodes_h_l2123_c7_7514_return_output,
 CONST_SR_8_uxn_opcodes_h_l2128_c31_d706_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2111_c3_2b7a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2106_c2_563f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2115_c3_c732 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2114_c7_4abc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2114_c7_4abc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2123_c7_7514_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2117_c7_d69f_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2123_c7_7514_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l2128_c31_d706_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l2128_c31_d706_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2128_c21_a728_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l2131_c3_5df4 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_return_output : unsigned(16 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2132_c21_5d31_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_d3c4_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_75a9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2117_l2106_l2114_DUPLICATE_3e64_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2106_l2123_l2114_DUPLICATE_77b0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2117_l2114_l2106_l2134_l2130_DUPLICATE_3d60_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2117_l2114_l2134_l2130_l2123_DUPLICATE_c3ac_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2117_l2114_DUPLICATE_2cef_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2_uxn_opcodes_h_l2139_l2102_DUPLICATE_0d85_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_right := to_unsigned(4, 3);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_y := to_signed(-4, 4);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_right := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2111_c3_2b7a := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2111_c3_2b7a;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2115_c3_c732 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2115_c3_c732;
     VAR_sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_right := to_unsigned(5, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_ins := VAR_ins;
     VAR_CONST_SR_8_uxn_opcodes_h_l2128_c31_d706_x := n16;
     VAR_n16_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_left := VAR_phase;
     VAR_n16_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue := VAR_previous_stack_read;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l2106_c6_ed3c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2117_l2114_l2106_l2134_l2130_DUPLICATE_3d60 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2117_l2114_l2106_l2134_l2130_DUPLICATE_3d60_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2130_c11_6548] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_left;
     BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_return_output := BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2134_c11_1b33] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_left;
     BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_return_output := BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_75a9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_75a9_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2106_l2123_l2114_DUPLICATE_77b0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2106_l2123_l2114_DUPLICATE_77b0_return_output := result.is_sp_shift;

     -- BIN_OP_PLUS[uxn_opcodes_h_l2131_c22_9913] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_left;
     BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_return_output := BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2121_c30_136a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_ins;
     sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_x;
     sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_return_output := sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2117_l2106_l2114_DUPLICATE_3e64 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2117_l2106_l2114_DUPLICATE_3e64_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2117_l2114_DUPLICATE_2cef LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2117_l2114_DUPLICATE_2cef_return_output := result.is_stack_operation_16bit;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2117_l2114_l2134_l2130_l2123_DUPLICATE_c3ac LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2117_l2114_l2134_l2130_l2123_DUPLICATE_c3ac_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2114_c11_f4ef] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_left;
     BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output := BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2117_c11_97d2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output;

     -- CONST_SR_8[uxn_opcodes_h_l2128_c31_d706] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l2128_c31_d706_x <= VAR_CONST_SR_8_uxn_opcodes_h_l2128_c31_d706_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l2128_c31_d706_return_output := CONST_SR_8_uxn_opcodes_h_l2128_c31_d706_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_d3c4 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_d3c4_return_output := result.u16_value;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2132_c21_5d31] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2132_c21_5d31_return_output := CAST_TO_uint8_t_uint16_t(
     n16);

     -- BIN_OP_EQ[uxn_opcodes_h_l2123_c11_18fe] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_left;
     BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_return_output := BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2114_c7_4abc] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2114_c7_4abc_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_n16_MUX_uxn_opcodes_h_l2106_c2_563f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2106_c2_563f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2106_c6_ed3c_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2114_c7_4abc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2114_c7_4abc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2114_c11_f4ef_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2117_c7_d69f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2117_c7_d69f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2117_c11_97d2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2123_c7_7514_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2123_c11_18fe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2130_c11_6548_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2134_c11_1b33_return_output;
     VAR_result_u16_value_uxn_opcodes_h_l2131_c3_5df4 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l2131_c22_9913_return_output, 16);
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2132_c21_5d31_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2117_l2106_l2114_DUPLICATE_3e64_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2117_l2106_l2114_DUPLICATE_3e64_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2117_l2106_l2114_DUPLICATE_3e64_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_d3c4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_d3c4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_d3c4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_d3c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2117_l2114_l2134_l2130_l2123_DUPLICATE_c3ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2117_l2114_l2134_l2130_l2123_DUPLICATE_c3ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2117_l2114_l2134_l2130_l2123_DUPLICATE_c3ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2117_l2114_l2134_l2130_l2123_DUPLICATE_c3ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2117_l2114_l2134_l2130_l2123_DUPLICATE_c3ac_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2117_l2114_l2106_l2134_l2130_DUPLICATE_3d60_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2117_l2114_l2106_l2134_l2130_DUPLICATE_3d60_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2117_l2114_l2106_l2134_l2130_DUPLICATE_3d60_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2117_l2114_l2106_l2134_l2130_DUPLICATE_3d60_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2117_l2114_l2106_l2134_l2130_DUPLICATE_3d60_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2106_l2123_l2114_DUPLICATE_77b0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2106_l2123_l2114_DUPLICATE_77b0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2106_l2123_l2114_DUPLICATE_77b0_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2117_l2114_DUPLICATE_2cef_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2117_l2114_DUPLICATE_2cef_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_75a9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_75a9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_75a9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2117_l2106_l2114_l2130_DUPLICATE_75a9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2114_c7_4abc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2121_c30_136a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue := VAR_result_u16_value_uxn_opcodes_h_l2131_c3_5df4;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2134_c7_a284] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2117_c7_d69f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2134_c7_a284] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2114_c7_4abc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2130_c7_333b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output := result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output;

     -- t16_MUX[uxn_opcodes_h_l2123_c7_7514] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2123_c7_7514_cond <= VAR_t16_MUX_uxn_opcodes_h_l2123_c7_7514_cond;
     t16_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue;
     t16_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2123_c7_7514_return_output := t16_MUX_uxn_opcodes_h_l2123_c7_7514_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2117_c7_d69f] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2130_c7_333b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2123_c7_7514] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2128_c21_a728] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2128_c21_a728_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l2128_c31_d706_return_output);

     -- n16_MUX[uxn_opcodes_h_l2117_c7_d69f] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2117_c7_d69f_cond <= VAR_n16_MUX_uxn_opcodes_h_l2117_c7_d69f_cond;
     n16_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue;
     n16_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output := n16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2128_c21_a728_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse := VAR_n16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2134_c7_a284_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2134_c7_a284_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2123_c7_7514_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2130_c7_333b_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2123_c7_7514_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2114_c7_4abc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2123_c7_7514] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output := result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2123_c7_7514] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output := result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2114_c7_4abc] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2106_c2_563f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2130_c7_333b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2117_c7_d69f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;

     -- n16_MUX[uxn_opcodes_h_l2114_c7_4abc] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2114_c7_4abc_cond <= VAR_n16_MUX_uxn_opcodes_h_l2114_c7_4abc_cond;
     n16_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue;
     n16_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output := n16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2130_c7_333b] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_return_output;

     -- t16_MUX[uxn_opcodes_h_l2117_c7_d69f] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2117_c7_d69f_cond <= VAR_t16_MUX_uxn_opcodes_h_l2117_c7_d69f_cond;
     t16_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue;
     t16_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output := t16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse := VAR_n16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2130_c7_333b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2130_c7_333b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2123_c7_7514_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2117_c7_d69f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2106_c2_563f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output;

     -- t16_MUX[uxn_opcodes_h_l2114_c7_4abc] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2114_c7_4abc_cond <= VAR_t16_MUX_uxn_opcodes_h_l2114_c7_4abc_cond;
     t16_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue;
     t16_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output := t16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2117_c7_d69f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output := result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2123_c7_7514] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_return_output;

     -- n16_MUX[uxn_opcodes_h_l2106_c2_563f] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2106_c2_563f_cond <= VAR_n16_MUX_uxn_opcodes_h_l2106_c2_563f_cond;
     n16_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue;
     n16_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output := n16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2114_c7_4abc] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2106_c2_563f] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2123_c7_7514] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_return_output;

     -- Submodule level 4
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2123_c7_7514_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2123_c7_7514_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l2114_c7_4abc] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output := result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2106_c2_563f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2114_c7_4abc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output := result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;

     -- t16_MUX[uxn_opcodes_h_l2106_c2_563f] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2106_c2_563f_cond <= VAR_t16_MUX_uxn_opcodes_h_l2106_c2_563f_cond;
     t16_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue;
     t16_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output := t16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2117_c7_d69f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2117_c7_d69f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2117_c7_d69f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2106_c2_563f_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l2106_c2_563f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output := result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2114_c7_4abc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2106_c2_563f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2114_c7_4abc] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2114_c7_4abc_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l2106_c2_563f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2106_c2_563f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2_uxn_opcodes_h_l2139_l2102_DUPLICATE_0d85 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2_uxn_opcodes_h_l2139_l2102_DUPLICATE_0d85_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2106_c2_563f_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2106_c2_563f_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2_uxn_opcodes_h_l2139_l2102_DUPLICATE_0d85_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2_uxn_opcodes_h_l2139_l2102_DUPLICATE_0d85_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
