-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 19
entity uint16_mux16_0CLK_4e6656cf is
port(
 sel : in unsigned(3 downto 0);
 in0 : in unsigned(15 downto 0);
 in1 : in unsigned(15 downto 0);
 in2 : in unsigned(15 downto 0);
 in3 : in unsigned(15 downto 0);
 in4 : in unsigned(15 downto 0);
 in5 : in unsigned(15 downto 0);
 in6 : in unsigned(15 downto 0);
 in7 : in unsigned(15 downto 0);
 in8 : in unsigned(15 downto 0);
 in9 : in unsigned(15 downto 0);
 in10 : in unsigned(15 downto 0);
 in11 : in unsigned(15 downto 0);
 in12 : in unsigned(15 downto 0);
 in13 : in unsigned(15 downto 0);
 in14 : in unsigned(15 downto 0);
 in15 : in unsigned(15 downto 0);
 return_output : out unsigned(15 downto 0));
end uint16_mux16_0CLK_4e6656cf;
architecture arch of uint16_mux16_0CLK_4e6656cf is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- layer0_node0_MUX[bit_math_h_l18_c3_07cc]
signal layer0_node0_MUX_bit_math_h_l18_c3_07cc_cond : unsigned(0 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_07cc_iftrue : unsigned(15 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_07cc_iffalse : unsigned(15 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_07cc_return_output : unsigned(15 downto 0);

-- layer0_node1_MUX[bit_math_h_l29_c3_bb0c]
signal layer0_node1_MUX_bit_math_h_l29_c3_bb0c_cond : unsigned(0 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_bb0c_iftrue : unsigned(15 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_bb0c_iffalse : unsigned(15 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_bb0c_return_output : unsigned(15 downto 0);

-- layer0_node2_MUX[bit_math_h_l40_c3_d671]
signal layer0_node2_MUX_bit_math_h_l40_c3_d671_cond : unsigned(0 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_d671_iftrue : unsigned(15 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_d671_iffalse : unsigned(15 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_d671_return_output : unsigned(15 downto 0);

-- layer0_node3_MUX[bit_math_h_l51_c3_0e8e]
signal layer0_node3_MUX_bit_math_h_l51_c3_0e8e_cond : unsigned(0 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_0e8e_iftrue : unsigned(15 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_0e8e_iffalse : unsigned(15 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_0e8e_return_output : unsigned(15 downto 0);

-- layer0_node4_MUX[bit_math_h_l62_c3_afa9]
signal layer0_node4_MUX_bit_math_h_l62_c3_afa9_cond : unsigned(0 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_afa9_iftrue : unsigned(15 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_afa9_iffalse : unsigned(15 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_afa9_return_output : unsigned(15 downto 0);

-- layer0_node5_MUX[bit_math_h_l73_c3_fc87]
signal layer0_node5_MUX_bit_math_h_l73_c3_fc87_cond : unsigned(0 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_fc87_iftrue : unsigned(15 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_fc87_iffalse : unsigned(15 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_fc87_return_output : unsigned(15 downto 0);

-- layer0_node6_MUX[bit_math_h_l84_c3_48cb]
signal layer0_node6_MUX_bit_math_h_l84_c3_48cb_cond : unsigned(0 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_48cb_iftrue : unsigned(15 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_48cb_iffalse : unsigned(15 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_48cb_return_output : unsigned(15 downto 0);

-- layer0_node7_MUX[bit_math_h_l95_c3_c04f]
signal layer0_node7_MUX_bit_math_h_l95_c3_c04f_cond : unsigned(0 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_c04f_iftrue : unsigned(15 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_c04f_iffalse : unsigned(15 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_c04f_return_output : unsigned(15 downto 0);

-- layer1_node0_MUX[bit_math_h_l112_c3_4341]
signal layer1_node0_MUX_bit_math_h_l112_c3_4341_cond : unsigned(0 downto 0);
signal layer1_node0_MUX_bit_math_h_l112_c3_4341_iftrue : unsigned(15 downto 0);
signal layer1_node0_MUX_bit_math_h_l112_c3_4341_iffalse : unsigned(15 downto 0);
signal layer1_node0_MUX_bit_math_h_l112_c3_4341_return_output : unsigned(15 downto 0);

-- layer1_node1_MUX[bit_math_h_l123_c3_88dc]
signal layer1_node1_MUX_bit_math_h_l123_c3_88dc_cond : unsigned(0 downto 0);
signal layer1_node1_MUX_bit_math_h_l123_c3_88dc_iftrue : unsigned(15 downto 0);
signal layer1_node1_MUX_bit_math_h_l123_c3_88dc_iffalse : unsigned(15 downto 0);
signal layer1_node1_MUX_bit_math_h_l123_c3_88dc_return_output : unsigned(15 downto 0);

-- layer1_node2_MUX[bit_math_h_l134_c3_ee56]
signal layer1_node2_MUX_bit_math_h_l134_c3_ee56_cond : unsigned(0 downto 0);
signal layer1_node2_MUX_bit_math_h_l134_c3_ee56_iftrue : unsigned(15 downto 0);
signal layer1_node2_MUX_bit_math_h_l134_c3_ee56_iffalse : unsigned(15 downto 0);
signal layer1_node2_MUX_bit_math_h_l134_c3_ee56_return_output : unsigned(15 downto 0);

-- layer1_node3_MUX[bit_math_h_l145_c3_2d21]
signal layer1_node3_MUX_bit_math_h_l145_c3_2d21_cond : unsigned(0 downto 0);
signal layer1_node3_MUX_bit_math_h_l145_c3_2d21_iftrue : unsigned(15 downto 0);
signal layer1_node3_MUX_bit_math_h_l145_c3_2d21_iffalse : unsigned(15 downto 0);
signal layer1_node3_MUX_bit_math_h_l145_c3_2d21_return_output : unsigned(15 downto 0);

-- layer2_node0_MUX[bit_math_h_l162_c3_ff65]
signal layer2_node0_MUX_bit_math_h_l162_c3_ff65_cond : unsigned(0 downto 0);
signal layer2_node0_MUX_bit_math_h_l162_c3_ff65_iftrue : unsigned(15 downto 0);
signal layer2_node0_MUX_bit_math_h_l162_c3_ff65_iffalse : unsigned(15 downto 0);
signal layer2_node0_MUX_bit_math_h_l162_c3_ff65_return_output : unsigned(15 downto 0);

-- layer2_node1_MUX[bit_math_h_l173_c3_2b00]
signal layer2_node1_MUX_bit_math_h_l173_c3_2b00_cond : unsigned(0 downto 0);
signal layer2_node1_MUX_bit_math_h_l173_c3_2b00_iftrue : unsigned(15 downto 0);
signal layer2_node1_MUX_bit_math_h_l173_c3_2b00_iffalse : unsigned(15 downto 0);
signal layer2_node1_MUX_bit_math_h_l173_c3_2b00_return_output : unsigned(15 downto 0);

-- layer3_node0_MUX[bit_math_h_l190_c3_ddd7]
signal layer3_node0_MUX_bit_math_h_l190_c3_ddd7_cond : unsigned(0 downto 0);
signal layer3_node0_MUX_bit_math_h_l190_c3_ddd7_iftrue : unsigned(15 downto 0);
signal layer3_node0_MUX_bit_math_h_l190_c3_ddd7_iffalse : unsigned(15 downto 0);
signal layer3_node0_MUX_bit_math_h_l190_c3_ddd7_return_output : unsigned(15 downto 0);

function uint4_0_0( x : unsigned) return unsigned is
--variable x : unsigned(3 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(0- i);
      end loop;
return return_output;
end function;

function uint4_1_1( x : unsigned) return unsigned is
--variable x : unsigned(3 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(1- i);
      end loop;
return return_output;
end function;

function uint4_2_2( x : unsigned) return unsigned is
--variable x : unsigned(3 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(2- i);
      end loop;
return return_output;
end function;

function uint4_3_3( x : unsigned) return unsigned is
--variable x : unsigned(3 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(3- i);
      end loop;
return return_output;
end function;


begin

-- SUBMODULE INSTANCES 
-- layer0_node0_MUX_bit_math_h_l18_c3_07cc
layer0_node0_MUX_bit_math_h_l18_c3_07cc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node0_MUX_bit_math_h_l18_c3_07cc_cond,
layer0_node0_MUX_bit_math_h_l18_c3_07cc_iftrue,
layer0_node0_MUX_bit_math_h_l18_c3_07cc_iffalse,
layer0_node0_MUX_bit_math_h_l18_c3_07cc_return_output);

-- layer0_node1_MUX_bit_math_h_l29_c3_bb0c
layer0_node1_MUX_bit_math_h_l29_c3_bb0c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node1_MUX_bit_math_h_l29_c3_bb0c_cond,
layer0_node1_MUX_bit_math_h_l29_c3_bb0c_iftrue,
layer0_node1_MUX_bit_math_h_l29_c3_bb0c_iffalse,
layer0_node1_MUX_bit_math_h_l29_c3_bb0c_return_output);

-- layer0_node2_MUX_bit_math_h_l40_c3_d671
layer0_node2_MUX_bit_math_h_l40_c3_d671 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node2_MUX_bit_math_h_l40_c3_d671_cond,
layer0_node2_MUX_bit_math_h_l40_c3_d671_iftrue,
layer0_node2_MUX_bit_math_h_l40_c3_d671_iffalse,
layer0_node2_MUX_bit_math_h_l40_c3_d671_return_output);

-- layer0_node3_MUX_bit_math_h_l51_c3_0e8e
layer0_node3_MUX_bit_math_h_l51_c3_0e8e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node3_MUX_bit_math_h_l51_c3_0e8e_cond,
layer0_node3_MUX_bit_math_h_l51_c3_0e8e_iftrue,
layer0_node3_MUX_bit_math_h_l51_c3_0e8e_iffalse,
layer0_node3_MUX_bit_math_h_l51_c3_0e8e_return_output);

-- layer0_node4_MUX_bit_math_h_l62_c3_afa9
layer0_node4_MUX_bit_math_h_l62_c3_afa9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node4_MUX_bit_math_h_l62_c3_afa9_cond,
layer0_node4_MUX_bit_math_h_l62_c3_afa9_iftrue,
layer0_node4_MUX_bit_math_h_l62_c3_afa9_iffalse,
layer0_node4_MUX_bit_math_h_l62_c3_afa9_return_output);

-- layer0_node5_MUX_bit_math_h_l73_c3_fc87
layer0_node5_MUX_bit_math_h_l73_c3_fc87 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node5_MUX_bit_math_h_l73_c3_fc87_cond,
layer0_node5_MUX_bit_math_h_l73_c3_fc87_iftrue,
layer0_node5_MUX_bit_math_h_l73_c3_fc87_iffalse,
layer0_node5_MUX_bit_math_h_l73_c3_fc87_return_output);

-- layer0_node6_MUX_bit_math_h_l84_c3_48cb
layer0_node6_MUX_bit_math_h_l84_c3_48cb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node6_MUX_bit_math_h_l84_c3_48cb_cond,
layer0_node6_MUX_bit_math_h_l84_c3_48cb_iftrue,
layer0_node6_MUX_bit_math_h_l84_c3_48cb_iffalse,
layer0_node6_MUX_bit_math_h_l84_c3_48cb_return_output);

-- layer0_node7_MUX_bit_math_h_l95_c3_c04f
layer0_node7_MUX_bit_math_h_l95_c3_c04f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer0_node7_MUX_bit_math_h_l95_c3_c04f_cond,
layer0_node7_MUX_bit_math_h_l95_c3_c04f_iftrue,
layer0_node7_MUX_bit_math_h_l95_c3_c04f_iffalse,
layer0_node7_MUX_bit_math_h_l95_c3_c04f_return_output);

-- layer1_node0_MUX_bit_math_h_l112_c3_4341
layer1_node0_MUX_bit_math_h_l112_c3_4341 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer1_node0_MUX_bit_math_h_l112_c3_4341_cond,
layer1_node0_MUX_bit_math_h_l112_c3_4341_iftrue,
layer1_node0_MUX_bit_math_h_l112_c3_4341_iffalse,
layer1_node0_MUX_bit_math_h_l112_c3_4341_return_output);

-- layer1_node1_MUX_bit_math_h_l123_c3_88dc
layer1_node1_MUX_bit_math_h_l123_c3_88dc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer1_node1_MUX_bit_math_h_l123_c3_88dc_cond,
layer1_node1_MUX_bit_math_h_l123_c3_88dc_iftrue,
layer1_node1_MUX_bit_math_h_l123_c3_88dc_iffalse,
layer1_node1_MUX_bit_math_h_l123_c3_88dc_return_output);

-- layer1_node2_MUX_bit_math_h_l134_c3_ee56
layer1_node2_MUX_bit_math_h_l134_c3_ee56 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer1_node2_MUX_bit_math_h_l134_c3_ee56_cond,
layer1_node2_MUX_bit_math_h_l134_c3_ee56_iftrue,
layer1_node2_MUX_bit_math_h_l134_c3_ee56_iffalse,
layer1_node2_MUX_bit_math_h_l134_c3_ee56_return_output);

-- layer1_node3_MUX_bit_math_h_l145_c3_2d21
layer1_node3_MUX_bit_math_h_l145_c3_2d21 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer1_node3_MUX_bit_math_h_l145_c3_2d21_cond,
layer1_node3_MUX_bit_math_h_l145_c3_2d21_iftrue,
layer1_node3_MUX_bit_math_h_l145_c3_2d21_iffalse,
layer1_node3_MUX_bit_math_h_l145_c3_2d21_return_output);

-- layer2_node0_MUX_bit_math_h_l162_c3_ff65
layer2_node0_MUX_bit_math_h_l162_c3_ff65 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer2_node0_MUX_bit_math_h_l162_c3_ff65_cond,
layer2_node0_MUX_bit_math_h_l162_c3_ff65_iftrue,
layer2_node0_MUX_bit_math_h_l162_c3_ff65_iffalse,
layer2_node0_MUX_bit_math_h_l162_c3_ff65_return_output);

-- layer2_node1_MUX_bit_math_h_l173_c3_2b00
layer2_node1_MUX_bit_math_h_l173_c3_2b00 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer2_node1_MUX_bit_math_h_l173_c3_2b00_cond,
layer2_node1_MUX_bit_math_h_l173_c3_2b00_iftrue,
layer2_node1_MUX_bit_math_h_l173_c3_2b00_iffalse,
layer2_node1_MUX_bit_math_h_l173_c3_2b00_return_output);

-- layer3_node0_MUX_bit_math_h_l190_c3_ddd7
layer3_node0_MUX_bit_math_h_l190_c3_ddd7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
layer3_node0_MUX_bit_math_h_l190_c3_ddd7_cond,
layer3_node0_MUX_bit_math_h_l190_c3_ddd7_iftrue,
layer3_node0_MUX_bit_math_h_l190_c3_ddd7_iffalse,
layer3_node0_MUX_bit_math_h_l190_c3_ddd7_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 sel,
 in0,
 in1,
 in2,
 in3,
 in4,
 in5,
 in6,
 in7,
 in8,
 in9,
 in10,
 in11,
 in12,
 in13,
 in14,
 in15,
 -- All submodule outputs
 layer0_node0_MUX_bit_math_h_l18_c3_07cc_return_output,
 layer0_node1_MUX_bit_math_h_l29_c3_bb0c_return_output,
 layer0_node2_MUX_bit_math_h_l40_c3_d671_return_output,
 layer0_node3_MUX_bit_math_h_l51_c3_0e8e_return_output,
 layer0_node4_MUX_bit_math_h_l62_c3_afa9_return_output,
 layer0_node5_MUX_bit_math_h_l73_c3_fc87_return_output,
 layer0_node6_MUX_bit_math_h_l84_c3_48cb_return_output,
 layer0_node7_MUX_bit_math_h_l95_c3_c04f_return_output,
 layer1_node0_MUX_bit_math_h_l112_c3_4341_return_output,
 layer1_node1_MUX_bit_math_h_l123_c3_88dc_return_output,
 layer1_node2_MUX_bit_math_h_l134_c3_ee56_return_output,
 layer1_node3_MUX_bit_math_h_l145_c3_2d21_return_output,
 layer2_node0_MUX_bit_math_h_l162_c3_ff65_return_output,
 layer2_node1_MUX_bit_math_h_l173_c3_2b00_return_output,
 layer3_node0_MUX_bit_math_h_l190_c3_ddd7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(15 downto 0);
 variable VAR_sel : unsigned(3 downto 0);
 variable VAR_in0 : unsigned(15 downto 0);
 variable VAR_in1 : unsigned(15 downto 0);
 variable VAR_in2 : unsigned(15 downto 0);
 variable VAR_in3 : unsigned(15 downto 0);
 variable VAR_in4 : unsigned(15 downto 0);
 variable VAR_in5 : unsigned(15 downto 0);
 variable VAR_in6 : unsigned(15 downto 0);
 variable VAR_in7 : unsigned(15 downto 0);
 variable VAR_in8 : unsigned(15 downto 0);
 variable VAR_in9 : unsigned(15 downto 0);
 variable VAR_in10 : unsigned(15 downto 0);
 variable VAR_in11 : unsigned(15 downto 0);
 variable VAR_in12 : unsigned(15 downto 0);
 variable VAR_in13 : unsigned(15 downto 0);
 variable VAR_in14 : unsigned(15 downto 0);
 variable VAR_in15 : unsigned(15 downto 0);
 variable VAR_sel0 : unsigned(0 downto 0);
 variable VAR_uint4_0_0_bit_math_h_l14_c10_7a75_return_output : unsigned(0 downto 0);
 variable VAR_layer0_node0 : unsigned(15 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_07cc_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_07cc_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_07cc_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_07cc_cond : unsigned(0 downto 0);
 variable VAR_layer0_node1 : unsigned(15 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_bb0c_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_bb0c_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_bb0c_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_bb0c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node2 : unsigned(15 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_d671_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_d671_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_d671_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_d671_cond : unsigned(0 downto 0);
 variable VAR_layer0_node3 : unsigned(15 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_0e8e_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_0e8e_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_0e8e_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_0e8e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node4 : unsigned(15 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_afa9_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_afa9_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_afa9_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_afa9_cond : unsigned(0 downto 0);
 variable VAR_layer0_node5 : unsigned(15 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_fc87_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_fc87_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_fc87_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_fc87_cond : unsigned(0 downto 0);
 variable VAR_layer0_node6 : unsigned(15 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_48cb_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_48cb_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_48cb_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_48cb_cond : unsigned(0 downto 0);
 variable VAR_layer0_node7 : unsigned(15 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_c04f_iftrue : unsigned(15 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_c04f_iffalse : unsigned(15 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_c04f_return_output : unsigned(15 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_c04f_cond : unsigned(0 downto 0);
 variable VAR_sel1 : unsigned(0 downto 0);
 variable VAR_uint4_1_1_bit_math_h_l108_c10_67d7_return_output : unsigned(0 downto 0);
 variable VAR_layer1_node0 : unsigned(15 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l112_c3_4341_iftrue : unsigned(15 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l112_c3_4341_iffalse : unsigned(15 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l112_c3_4341_return_output : unsigned(15 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l112_c3_4341_cond : unsigned(0 downto 0);
 variable VAR_layer1_node1 : unsigned(15 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l123_c3_88dc_iftrue : unsigned(15 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l123_c3_88dc_iffalse : unsigned(15 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l123_c3_88dc_return_output : unsigned(15 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l123_c3_88dc_cond : unsigned(0 downto 0);
 variable VAR_layer1_node2 : unsigned(15 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l134_c3_ee56_iftrue : unsigned(15 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l134_c3_ee56_iffalse : unsigned(15 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l134_c3_ee56_return_output : unsigned(15 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l134_c3_ee56_cond : unsigned(0 downto 0);
 variable VAR_layer1_node3 : unsigned(15 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l145_c3_2d21_iftrue : unsigned(15 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l145_c3_2d21_iffalse : unsigned(15 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l145_c3_2d21_return_output : unsigned(15 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l145_c3_2d21_cond : unsigned(0 downto 0);
 variable VAR_sel2 : unsigned(0 downto 0);
 variable VAR_uint4_2_2_bit_math_h_l158_c10_bf6d_return_output : unsigned(0 downto 0);
 variable VAR_layer2_node0 : unsigned(15 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l162_c3_ff65_iftrue : unsigned(15 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l162_c3_ff65_iffalse : unsigned(15 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l162_c3_ff65_return_output : unsigned(15 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l162_c3_ff65_cond : unsigned(0 downto 0);
 variable VAR_layer2_node1 : unsigned(15 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l173_c3_2b00_iftrue : unsigned(15 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l173_c3_2b00_iffalse : unsigned(15 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l173_c3_2b00_return_output : unsigned(15 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l173_c3_2b00_cond : unsigned(0 downto 0);
 variable VAR_sel3 : unsigned(0 downto 0);
 variable VAR_uint4_3_3_bit_math_h_l186_c10_017f_return_output : unsigned(0 downto 0);
 variable VAR_layer3_node0 : unsigned(15 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l190_c3_ddd7_iftrue : unsigned(15 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l190_c3_ddd7_iffalse : unsigned(15 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l190_c3_ddd7_return_output : unsigned(15 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l190_c3_ddd7_cond : unsigned(0 downto 0);
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_sel := sel;
     VAR_in0 := in0;
     VAR_in1 := in1;
     VAR_in2 := in2;
     VAR_in3 := in3;
     VAR_in4 := in4;
     VAR_in5 := in5;
     VAR_in6 := in6;
     VAR_in7 := in7;
     VAR_in8 := in8;
     VAR_in9 := in9;
     VAR_in10 := in10;
     VAR_in11 := in11;
     VAR_in12 := in12;
     VAR_in13 := in13;
     VAR_in14 := in14;
     VAR_in15 := in15;

     -- Submodule level 0
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_07cc_iffalse := VAR_in0;
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_07cc_iftrue := VAR_in1;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_fc87_iffalse := VAR_in10;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_fc87_iftrue := VAR_in11;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_48cb_iffalse := VAR_in12;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_48cb_iftrue := VAR_in13;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_c04f_iffalse := VAR_in14;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_c04f_iftrue := VAR_in15;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_bb0c_iffalse := VAR_in2;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_bb0c_iftrue := VAR_in3;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_d671_iffalse := VAR_in4;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_d671_iftrue := VAR_in5;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_0e8e_iffalse := VAR_in6;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_0e8e_iftrue := VAR_in7;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_afa9_iffalse := VAR_in8;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_afa9_iftrue := VAR_in9;
     -- uint4_0_0[bit_math_h_l14_c10_7a75] LATENCY=0
     VAR_uint4_0_0_bit_math_h_l14_c10_7a75_return_output := uint4_0_0(
     VAR_sel);

     -- uint4_3_3[bit_math_h_l186_c10_017f] LATENCY=0
     VAR_uint4_3_3_bit_math_h_l186_c10_017f_return_output := uint4_3_3(
     VAR_sel);

     -- uint4_1_1[bit_math_h_l108_c10_67d7] LATENCY=0
     VAR_uint4_1_1_bit_math_h_l108_c10_67d7_return_output := uint4_1_1(
     VAR_sel);

     -- uint4_2_2[bit_math_h_l158_c10_bf6d] LATENCY=0
     VAR_uint4_2_2_bit_math_h_l158_c10_bf6d_return_output := uint4_2_2(
     VAR_sel);

     -- Submodule level 1
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_07cc_cond := VAR_uint4_0_0_bit_math_h_l14_c10_7a75_return_output;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_bb0c_cond := VAR_uint4_0_0_bit_math_h_l14_c10_7a75_return_output;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_d671_cond := VAR_uint4_0_0_bit_math_h_l14_c10_7a75_return_output;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_0e8e_cond := VAR_uint4_0_0_bit_math_h_l14_c10_7a75_return_output;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_afa9_cond := VAR_uint4_0_0_bit_math_h_l14_c10_7a75_return_output;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_fc87_cond := VAR_uint4_0_0_bit_math_h_l14_c10_7a75_return_output;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_48cb_cond := VAR_uint4_0_0_bit_math_h_l14_c10_7a75_return_output;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_c04f_cond := VAR_uint4_0_0_bit_math_h_l14_c10_7a75_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l112_c3_4341_cond := VAR_uint4_1_1_bit_math_h_l108_c10_67d7_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l123_c3_88dc_cond := VAR_uint4_1_1_bit_math_h_l108_c10_67d7_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l134_c3_ee56_cond := VAR_uint4_1_1_bit_math_h_l108_c10_67d7_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l145_c3_2d21_cond := VAR_uint4_1_1_bit_math_h_l108_c10_67d7_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l162_c3_ff65_cond := VAR_uint4_2_2_bit_math_h_l158_c10_bf6d_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l173_c3_2b00_cond := VAR_uint4_2_2_bit_math_h_l158_c10_bf6d_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l190_c3_ddd7_cond := VAR_uint4_3_3_bit_math_h_l186_c10_017f_return_output;
     -- layer0_node6_MUX[bit_math_h_l84_c3_48cb] LATENCY=0
     -- Inputs
     layer0_node6_MUX_bit_math_h_l84_c3_48cb_cond <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_48cb_cond;
     layer0_node6_MUX_bit_math_h_l84_c3_48cb_iftrue <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_48cb_iftrue;
     layer0_node6_MUX_bit_math_h_l84_c3_48cb_iffalse <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_48cb_iffalse;
     -- Outputs
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_48cb_return_output := layer0_node6_MUX_bit_math_h_l84_c3_48cb_return_output;

     -- layer0_node7_MUX[bit_math_h_l95_c3_c04f] LATENCY=0
     -- Inputs
     layer0_node7_MUX_bit_math_h_l95_c3_c04f_cond <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_c04f_cond;
     layer0_node7_MUX_bit_math_h_l95_c3_c04f_iftrue <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_c04f_iftrue;
     layer0_node7_MUX_bit_math_h_l95_c3_c04f_iffalse <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_c04f_iffalse;
     -- Outputs
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_c04f_return_output := layer0_node7_MUX_bit_math_h_l95_c3_c04f_return_output;

     -- layer0_node5_MUX[bit_math_h_l73_c3_fc87] LATENCY=0
     -- Inputs
     layer0_node5_MUX_bit_math_h_l73_c3_fc87_cond <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_fc87_cond;
     layer0_node5_MUX_bit_math_h_l73_c3_fc87_iftrue <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_fc87_iftrue;
     layer0_node5_MUX_bit_math_h_l73_c3_fc87_iffalse <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_fc87_iffalse;
     -- Outputs
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_fc87_return_output := layer0_node5_MUX_bit_math_h_l73_c3_fc87_return_output;

     -- layer0_node0_MUX[bit_math_h_l18_c3_07cc] LATENCY=0
     -- Inputs
     layer0_node0_MUX_bit_math_h_l18_c3_07cc_cond <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_07cc_cond;
     layer0_node0_MUX_bit_math_h_l18_c3_07cc_iftrue <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_07cc_iftrue;
     layer0_node0_MUX_bit_math_h_l18_c3_07cc_iffalse <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_07cc_iffalse;
     -- Outputs
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_07cc_return_output := layer0_node0_MUX_bit_math_h_l18_c3_07cc_return_output;

     -- layer0_node3_MUX[bit_math_h_l51_c3_0e8e] LATENCY=0
     -- Inputs
     layer0_node3_MUX_bit_math_h_l51_c3_0e8e_cond <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_0e8e_cond;
     layer0_node3_MUX_bit_math_h_l51_c3_0e8e_iftrue <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_0e8e_iftrue;
     layer0_node3_MUX_bit_math_h_l51_c3_0e8e_iffalse <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_0e8e_iffalse;
     -- Outputs
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_0e8e_return_output := layer0_node3_MUX_bit_math_h_l51_c3_0e8e_return_output;

     -- layer0_node2_MUX[bit_math_h_l40_c3_d671] LATENCY=0
     -- Inputs
     layer0_node2_MUX_bit_math_h_l40_c3_d671_cond <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_d671_cond;
     layer0_node2_MUX_bit_math_h_l40_c3_d671_iftrue <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_d671_iftrue;
     layer0_node2_MUX_bit_math_h_l40_c3_d671_iffalse <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_d671_iffalse;
     -- Outputs
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_d671_return_output := layer0_node2_MUX_bit_math_h_l40_c3_d671_return_output;

     -- layer0_node1_MUX[bit_math_h_l29_c3_bb0c] LATENCY=0
     -- Inputs
     layer0_node1_MUX_bit_math_h_l29_c3_bb0c_cond <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_bb0c_cond;
     layer0_node1_MUX_bit_math_h_l29_c3_bb0c_iftrue <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_bb0c_iftrue;
     layer0_node1_MUX_bit_math_h_l29_c3_bb0c_iffalse <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_bb0c_iffalse;
     -- Outputs
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_bb0c_return_output := layer0_node1_MUX_bit_math_h_l29_c3_bb0c_return_output;

     -- layer0_node4_MUX[bit_math_h_l62_c3_afa9] LATENCY=0
     -- Inputs
     layer0_node4_MUX_bit_math_h_l62_c3_afa9_cond <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_afa9_cond;
     layer0_node4_MUX_bit_math_h_l62_c3_afa9_iftrue <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_afa9_iftrue;
     layer0_node4_MUX_bit_math_h_l62_c3_afa9_iffalse <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_afa9_iffalse;
     -- Outputs
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_afa9_return_output := layer0_node4_MUX_bit_math_h_l62_c3_afa9_return_output;

     -- Submodule level 2
     VAR_layer1_node0_MUX_bit_math_h_l112_c3_4341_iffalse := VAR_layer0_node0_MUX_bit_math_h_l18_c3_07cc_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l112_c3_4341_iftrue := VAR_layer0_node1_MUX_bit_math_h_l29_c3_bb0c_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l123_c3_88dc_iffalse := VAR_layer0_node2_MUX_bit_math_h_l40_c3_d671_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l123_c3_88dc_iftrue := VAR_layer0_node3_MUX_bit_math_h_l51_c3_0e8e_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l134_c3_ee56_iffalse := VAR_layer0_node4_MUX_bit_math_h_l62_c3_afa9_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l134_c3_ee56_iftrue := VAR_layer0_node5_MUX_bit_math_h_l73_c3_fc87_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l145_c3_2d21_iffalse := VAR_layer0_node6_MUX_bit_math_h_l84_c3_48cb_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l145_c3_2d21_iftrue := VAR_layer0_node7_MUX_bit_math_h_l95_c3_c04f_return_output;
     -- layer1_node2_MUX[bit_math_h_l134_c3_ee56] LATENCY=0
     -- Inputs
     layer1_node2_MUX_bit_math_h_l134_c3_ee56_cond <= VAR_layer1_node2_MUX_bit_math_h_l134_c3_ee56_cond;
     layer1_node2_MUX_bit_math_h_l134_c3_ee56_iftrue <= VAR_layer1_node2_MUX_bit_math_h_l134_c3_ee56_iftrue;
     layer1_node2_MUX_bit_math_h_l134_c3_ee56_iffalse <= VAR_layer1_node2_MUX_bit_math_h_l134_c3_ee56_iffalse;
     -- Outputs
     VAR_layer1_node2_MUX_bit_math_h_l134_c3_ee56_return_output := layer1_node2_MUX_bit_math_h_l134_c3_ee56_return_output;

     -- layer1_node0_MUX[bit_math_h_l112_c3_4341] LATENCY=0
     -- Inputs
     layer1_node0_MUX_bit_math_h_l112_c3_4341_cond <= VAR_layer1_node0_MUX_bit_math_h_l112_c3_4341_cond;
     layer1_node0_MUX_bit_math_h_l112_c3_4341_iftrue <= VAR_layer1_node0_MUX_bit_math_h_l112_c3_4341_iftrue;
     layer1_node0_MUX_bit_math_h_l112_c3_4341_iffalse <= VAR_layer1_node0_MUX_bit_math_h_l112_c3_4341_iffalse;
     -- Outputs
     VAR_layer1_node0_MUX_bit_math_h_l112_c3_4341_return_output := layer1_node0_MUX_bit_math_h_l112_c3_4341_return_output;

     -- layer1_node1_MUX[bit_math_h_l123_c3_88dc] LATENCY=0
     -- Inputs
     layer1_node1_MUX_bit_math_h_l123_c3_88dc_cond <= VAR_layer1_node1_MUX_bit_math_h_l123_c3_88dc_cond;
     layer1_node1_MUX_bit_math_h_l123_c3_88dc_iftrue <= VAR_layer1_node1_MUX_bit_math_h_l123_c3_88dc_iftrue;
     layer1_node1_MUX_bit_math_h_l123_c3_88dc_iffalse <= VAR_layer1_node1_MUX_bit_math_h_l123_c3_88dc_iffalse;
     -- Outputs
     VAR_layer1_node1_MUX_bit_math_h_l123_c3_88dc_return_output := layer1_node1_MUX_bit_math_h_l123_c3_88dc_return_output;

     -- layer1_node3_MUX[bit_math_h_l145_c3_2d21] LATENCY=0
     -- Inputs
     layer1_node3_MUX_bit_math_h_l145_c3_2d21_cond <= VAR_layer1_node3_MUX_bit_math_h_l145_c3_2d21_cond;
     layer1_node3_MUX_bit_math_h_l145_c3_2d21_iftrue <= VAR_layer1_node3_MUX_bit_math_h_l145_c3_2d21_iftrue;
     layer1_node3_MUX_bit_math_h_l145_c3_2d21_iffalse <= VAR_layer1_node3_MUX_bit_math_h_l145_c3_2d21_iffalse;
     -- Outputs
     VAR_layer1_node3_MUX_bit_math_h_l145_c3_2d21_return_output := layer1_node3_MUX_bit_math_h_l145_c3_2d21_return_output;

     -- Submodule level 3
     VAR_layer2_node0_MUX_bit_math_h_l162_c3_ff65_iffalse := VAR_layer1_node0_MUX_bit_math_h_l112_c3_4341_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l162_c3_ff65_iftrue := VAR_layer1_node1_MUX_bit_math_h_l123_c3_88dc_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l173_c3_2b00_iffalse := VAR_layer1_node2_MUX_bit_math_h_l134_c3_ee56_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l173_c3_2b00_iftrue := VAR_layer1_node3_MUX_bit_math_h_l145_c3_2d21_return_output;
     -- layer2_node1_MUX[bit_math_h_l173_c3_2b00] LATENCY=0
     -- Inputs
     layer2_node1_MUX_bit_math_h_l173_c3_2b00_cond <= VAR_layer2_node1_MUX_bit_math_h_l173_c3_2b00_cond;
     layer2_node1_MUX_bit_math_h_l173_c3_2b00_iftrue <= VAR_layer2_node1_MUX_bit_math_h_l173_c3_2b00_iftrue;
     layer2_node1_MUX_bit_math_h_l173_c3_2b00_iffalse <= VAR_layer2_node1_MUX_bit_math_h_l173_c3_2b00_iffalse;
     -- Outputs
     VAR_layer2_node1_MUX_bit_math_h_l173_c3_2b00_return_output := layer2_node1_MUX_bit_math_h_l173_c3_2b00_return_output;

     -- layer2_node0_MUX[bit_math_h_l162_c3_ff65] LATENCY=0
     -- Inputs
     layer2_node0_MUX_bit_math_h_l162_c3_ff65_cond <= VAR_layer2_node0_MUX_bit_math_h_l162_c3_ff65_cond;
     layer2_node0_MUX_bit_math_h_l162_c3_ff65_iftrue <= VAR_layer2_node0_MUX_bit_math_h_l162_c3_ff65_iftrue;
     layer2_node0_MUX_bit_math_h_l162_c3_ff65_iffalse <= VAR_layer2_node0_MUX_bit_math_h_l162_c3_ff65_iffalse;
     -- Outputs
     VAR_layer2_node0_MUX_bit_math_h_l162_c3_ff65_return_output := layer2_node0_MUX_bit_math_h_l162_c3_ff65_return_output;

     -- Submodule level 4
     VAR_layer3_node0_MUX_bit_math_h_l190_c3_ddd7_iffalse := VAR_layer2_node0_MUX_bit_math_h_l162_c3_ff65_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l190_c3_ddd7_iftrue := VAR_layer2_node1_MUX_bit_math_h_l173_c3_2b00_return_output;
     -- layer3_node0_MUX[bit_math_h_l190_c3_ddd7] LATENCY=0
     -- Inputs
     layer3_node0_MUX_bit_math_h_l190_c3_ddd7_cond <= VAR_layer3_node0_MUX_bit_math_h_l190_c3_ddd7_cond;
     layer3_node0_MUX_bit_math_h_l190_c3_ddd7_iftrue <= VAR_layer3_node0_MUX_bit_math_h_l190_c3_ddd7_iftrue;
     layer3_node0_MUX_bit_math_h_l190_c3_ddd7_iffalse <= VAR_layer3_node0_MUX_bit_math_h_l190_c3_ddd7_iffalse;
     -- Outputs
     VAR_layer3_node0_MUX_bit_math_h_l190_c3_ddd7_return_output := layer3_node0_MUX_bit_math_h_l190_c3_ddd7_return_output;

     -- Submodule level 5
     VAR_return_output := VAR_layer3_node0_MUX_bit_math_h_l190_c3_ddd7_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
