-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 33
entity inc2_0CLK_d4b33a56 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end inc2_0CLK_d4b33a56;
architecture arch of inc2_0CLK_d4b33a56 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1228_c6_5d9d]
signal BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1228_c2_9878]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1228_c2_9878]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1228_c2_9878]
signal result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1228_c2_9878]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1228_c2_9878]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1228_c2_9878]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1228_c2_9878]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l1228_c2_9878]
signal t16_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1236_c11_2255]
signal BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1236_c7_a040]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1236_c7_a040]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1236_c7_a040]
signal result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1236_c7_a040]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1236_c7_a040]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1236_c7_a040]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1236_c7_a040]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l1236_c7_a040]
signal t16_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1238_c30_fb6e]
signal sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1240_c11_e4ae]
signal BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1240_c7_88ae]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1240_c7_88ae]
signal result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1240_c7_88ae]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1240_c7_88ae]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1240_c7_88ae]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1240_c7_88ae]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(3 downto 0);

-- t16_MUX[uxn_opcodes_h_l1240_c7_88ae]
signal t16_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1245_c22_bde3]
signal BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1247_c11_8f80]
signal BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1247_c7_91d9]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1247_c7_91d9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1247_c7_91d9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d
BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_left,
BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_right,
BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878
result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878
result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_cond,
result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878
result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878
result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878
result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_return_output);

-- t16_MUX_uxn_opcodes_h_l1228_c2_9878
t16_MUX_uxn_opcodes_h_l1228_c2_9878 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1228_c2_9878_cond,
t16_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue,
t16_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse,
t16_MUX_uxn_opcodes_h_l1228_c2_9878_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255
BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_left,
BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_right,
BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040
result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040
result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_cond,
result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040
result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040
result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040
result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_return_output);

-- t16_MUX_uxn_opcodes_h_l1236_c7_a040
t16_MUX_uxn_opcodes_h_l1236_c7_a040 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1236_c7_a040_cond,
t16_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue,
t16_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse,
t16_MUX_uxn_opcodes_h_l1236_c7_a040_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e
sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_ins,
sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_x,
sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_y,
sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae
BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_left,
BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_right,
BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae
result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae
result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_cond,
result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae
result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae
result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output);

-- t16_MUX_uxn_opcodes_h_l1240_c7_88ae
t16_MUX_uxn_opcodes_h_l1240_c7_88ae : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1240_c7_88ae_cond,
t16_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue,
t16_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse,
t16_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3
BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3 : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_left,
BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_right,
BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80
BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_left,
BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_right,
BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9
result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9
result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
 t16_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_return_output,
 t16_MUX_uxn_opcodes_h_l1236_c7_a040_return_output,
 sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output,
 t16_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1232_c3_4eff : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1236_c7_a040_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1228_c2_9878_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1228_c2_9878_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1236_c7_a040_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1245_c3_2f80 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1244_c3_cec4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1240_c7_88ae_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1228_l1240_DUPLICATE_5608_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1228_l1240_l1236_DUPLICATE_f9ce_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1228_l1236_DUPLICATE_3ecb_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1228_l1247_l1236_DUPLICATE_d3f4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1240_l1236_DUPLICATE_3265_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1240_l1247_l1236_DUPLICATE_a614_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1240_l1247_l1236_DUPLICATE_1d0c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1253_l1224_DUPLICATE_a4db_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1232_c3_4eff := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1232_c3_4eff;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1244_c3_cec4 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1244_c3_cec4;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_right := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_left := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse := t16;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1228_l1236_DUPLICATE_3ecb LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1228_l1236_DUPLICATE_3ecb_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1240_l1247_l1236_DUPLICATE_1d0c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1240_l1247_l1236_DUPLICATE_1d0c_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1228_l1247_l1236_DUPLICATE_d3f4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1228_l1247_l1236_DUPLICATE_d3f4_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1247_c11_8f80] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_left;
     BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_return_output := BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1228_l1240_l1236_DUPLICATE_f9ce LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1228_l1240_l1236_DUPLICATE_f9ce_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1228_c6_5d9d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1240_c11_e4ae] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_left;
     BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_return_output := BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1240_l1247_l1236_DUPLICATE_a614 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1240_l1247_l1236_DUPLICATE_a614_return_output := result.is_stack_operation_16bit;

     -- BIN_OP_EQ[uxn_opcodes_h_l1236_c11_2255] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_left;
     BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output := BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1245_c22_bde3] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1238_c30_fb6e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_ins;
     sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_x;
     sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_return_output := sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1228_l1240_DUPLICATE_5608 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1228_l1240_DUPLICATE_5608_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1240_l1236_DUPLICATE_3265 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1240_l1236_DUPLICATE_3265_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1228_c2_9878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c6_5d9d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1236_c7_a040_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_2255_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1240_c7_88ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1240_c11_e4ae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1247_c11_8f80_return_output;
     VAR_result_u16_value_uxn_opcodes_h_l1245_c3_2f80 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1245_c22_bde3_return_output, 16);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1228_l1236_DUPLICATE_3ecb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1228_l1236_DUPLICATE_3ecb_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1228_l1240_l1236_DUPLICATE_f9ce_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1228_l1240_l1236_DUPLICATE_f9ce_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1228_l1240_l1236_DUPLICATE_f9ce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1240_l1247_l1236_DUPLICATE_1d0c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1240_l1247_l1236_DUPLICATE_1d0c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1240_l1247_l1236_DUPLICATE_1d0c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1228_l1240_DUPLICATE_5608_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1228_l1240_DUPLICATE_5608_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1240_l1247_l1236_DUPLICATE_a614_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1240_l1247_l1236_DUPLICATE_a614_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1240_l1247_l1236_DUPLICATE_a614_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1228_l1247_l1236_DUPLICATE_d3f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1228_l1247_l1236_DUPLICATE_d3f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1228_l1247_l1236_DUPLICATE_d3f4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1240_l1236_DUPLICATE_3265_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1240_l1236_DUPLICATE_3265_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1238_c30_fb6e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1245_c3_2f80;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1236_c7_a040] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1247_c7_91d9] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1240_c7_88ae] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1240_c7_88ae] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1247_c7_91d9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output;

     -- t16_MUX[uxn_opcodes_h_l1240_c7_88ae] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1240_c7_88ae_cond <= VAR_t16_MUX_uxn_opcodes_h_l1240_c7_88ae_cond;
     t16_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue;
     t16_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output := t16_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1240_c7_88ae] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output := result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1247_c7_91d9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1247_c7_91d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1236_c7_a040] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1240_c7_88ae] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;

     -- t16_MUX[uxn_opcodes_h_l1236_c7_a040] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1236_c7_a040_cond <= VAR_t16_MUX_uxn_opcodes_h_l1236_c7_a040_cond;
     t16_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue;
     t16_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1236_c7_a040_return_output := t16_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1228_c2_9878] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1240_c7_88ae] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1236_c7_a040] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_return_output := result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1236_c7_a040] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1240_c7_88ae] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1240_c7_88ae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1228_c2_9878] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_return_output := result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1228_c2_9878] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1236_c7_a040] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1236_c7_a040] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1228_c2_9878] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1236_c7_a040] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;

     -- t16_MUX[uxn_opcodes_h_l1228_c2_9878] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1228_c2_9878_cond <= VAR_t16_MUX_uxn_opcodes_h_l1228_c2_9878_cond;
     t16_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue;
     t16_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1228_c2_9878_return_output := t16_MUX_uxn_opcodes_h_l1228_c2_9878_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_a040_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l1228_c2_9878_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1228_c2_9878] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1228_c2_9878] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1228_c2_9878] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_return_output;

     -- Submodule level 5
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1253_l1224_DUPLICATE_a4db LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1253_l1224_DUPLICATE_a4db_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c2_9878_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c2_9878_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1253_l1224_DUPLICATE_a4db_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1253_l1224_DUPLICATE_a4db_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
