-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity div2_0CLK_4496d276 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end div2_0CLK_4496d276;
architecture arch of div2_0CLK_4496d276 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1896_c6_819b]
signal BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1896_c2_257d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1896_c2_257d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1896_c2_257d]
signal result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1896_c2_257d]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1896_c2_257d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1896_c2_257d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1896_c2_257d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1896_c2_257d]
signal n16_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1896_c2_257d]
signal tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1896_c2_257d]
signal t16_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1904_c11_d436]
signal BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1904_c7_e7dd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1904_c7_e7dd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1904_c7_e7dd]
signal result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1904_c7_e7dd]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1904_c7_e7dd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1904_c7_e7dd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1904_c7_e7dd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1904_c7_e7dd]
signal n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1904_c7_e7dd]
signal tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1904_c7_e7dd]
signal t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1907_c11_f74f]
signal BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1907_c7_71a7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1907_c7_71a7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1907_c7_71a7]
signal result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1907_c7_71a7]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1907_c7_71a7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1907_c7_71a7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1907_c7_71a7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1907_c7_71a7]
signal n16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1907_c7_71a7]
signal tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1907_c7_71a7]
signal t16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1910_c30_a0a9]
signal sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1912_c11_e71f]
signal BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1912_c7_bb1d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1912_c7_bb1d]
signal result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1912_c7_bb1d]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1912_c7_bb1d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1912_c7_bb1d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1912_c7_bb1d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l1912_c7_bb1d]
signal n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1912_c7_bb1d]
signal tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1914_c11_9bf3]
signal BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_left : unsigned(15 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_return_output : unsigned(0 downto 0);

-- BIN_OP_DIV[uxn_opcodes_h_l1914_c26_c14d]
signal BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_left : unsigned(15 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_right : unsigned(15 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_return_output : unsigned(15 downto 0);

-- MUX[uxn_opcodes_h_l1914_c11_ba09]
signal MUX_uxn_opcodes_h_l1914_c11_ba09_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1914_c11_ba09_iftrue : unsigned(15 downto 0);
signal MUX_uxn_opcodes_h_l1914_c11_ba09_iffalse : unsigned(15 downto 0);
signal MUX_uxn_opcodes_h_l1914_c11_ba09_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1920_c11_0923]
signal BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1920_c7_8e01]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1920_c7_8e01]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1920_c7_8e01]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b
BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_left,
BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_right,
BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d
result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d
result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_cond,
result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d
result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d
result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_return_output);

-- n16_MUX_uxn_opcodes_h_l1896_c2_257d
n16_MUX_uxn_opcodes_h_l1896_c2_257d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1896_c2_257d_cond,
n16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue,
n16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse,
n16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1896_c2_257d
tmp16_MUX_uxn_opcodes_h_l1896_c2_257d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_cond,
tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue,
tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse,
tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output);

-- t16_MUX_uxn_opcodes_h_l1896_c2_257d
t16_MUX_uxn_opcodes_h_l1896_c2_257d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1896_c2_257d_cond,
t16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue,
t16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse,
t16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436
BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_left,
BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_right,
BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd
result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd
result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond,
result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd
result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd
result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd
result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output);

-- n16_MUX_uxn_opcodes_h_l1904_c7_e7dd
n16_MUX_uxn_opcodes_h_l1904_c7_e7dd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond,
n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue,
n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse,
n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd
tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond,
tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue,
tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse,
tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output);

-- t16_MUX_uxn_opcodes_h_l1904_c7_e7dd
t16_MUX_uxn_opcodes_h_l1904_c7_e7dd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond,
t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue,
t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse,
t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f
BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_left,
BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_right,
BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7
result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7
result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_cond,
result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7
result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7
result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7
result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output);

-- n16_MUX_uxn_opcodes_h_l1907_c7_71a7
n16_MUX_uxn_opcodes_h_l1907_c7_71a7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond,
n16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue,
n16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse,
n16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7
tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond,
tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue,
tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse,
tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output);

-- t16_MUX_uxn_opcodes_h_l1907_c7_71a7
t16_MUX_uxn_opcodes_h_l1907_c7_71a7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond,
t16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue,
t16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse,
t16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9
sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_ins,
sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_x,
sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_y,
sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f
BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_left,
BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_right,
BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d
result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d
result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond,
result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output);

-- n16_MUX_uxn_opcodes_h_l1912_c7_bb1d
n16_MUX_uxn_opcodes_h_l1912_c7_bb1d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond,
n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue,
n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse,
n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d
tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond,
tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue,
tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse,
tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3
BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3 : entity work.BIN_OP_EQ_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_left,
BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_right,
BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_return_output);

-- BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d
BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d : entity work.BIN_OP_DIV_uint16_t_uint16_t_0CLK_2b0015ee port map (
BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_left,
BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_right,
BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_return_output);

-- MUX_uxn_opcodes_h_l1914_c11_ba09
MUX_uxn_opcodes_h_l1914_c11_ba09 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1914_c11_ba09_cond,
MUX_uxn_opcodes_h_l1914_c11_ba09_iftrue,
MUX_uxn_opcodes_h_l1914_c11_ba09_iffalse,
MUX_uxn_opcodes_h_l1914_c11_ba09_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923
BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_left,
BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_right,
BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01
result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01
result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
 n16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
 tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
 t16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output,
 n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output,
 tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output,
 t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output,
 n16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output,
 tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output,
 t16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output,
 sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output,
 n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output,
 tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_return_output,
 BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_return_output,
 MUX_uxn_opcodes_h_l1914_c11_ba09_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1901_c3_0b3b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1896_c2_257d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1905_c3_2d67 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1917_c3_e756 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1914_c11_ba09_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1914_c11_ba09_iftrue : unsigned(15 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1914_c11_ba09_iffalse : unsigned(15 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_return_output : unsigned(15 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1914_c11_ba09_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1912_l1904_l1896_DUPLICATE_abe2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1912_l1904_l1907_l1896_DUPLICATE_db41_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1904_l1907_l1896_DUPLICATE_68d6_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1904_l1920_l1907_l1896_DUPLICATE_0223_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_9571_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_398f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1912_l1907_DUPLICATE_a08c_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1926_l1892_DUPLICATE_8d40_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1905_c3_2d67 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1905_c3_2d67;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1917_c3_e756 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1917_c3_e756;
     VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_right := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1901_c3_0b3b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1901_c3_0b3b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_y := resize(to_signed(-2, 3), 4);
     VAR_MUX_uxn_opcodes_h_l1914_c11_ba09_iftrue := resize(to_unsigned(0, 1), 16);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_right := to_unsigned(4, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_left := VAR_phase;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_left := VAR_previous_stack_read;
     VAR_n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_right := t16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse := t16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse := tmp16;
     -- BIN_OP_EQ[uxn_opcodes_h_l1896_c6_819b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1904_c11_d436] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_left;
     BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output := BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1910_c30_a0a9] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_ins;
     sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_x;
     sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_return_output := sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1912_c11_e71f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1914_c11_9bf3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1912_l1904_l1907_l1896_DUPLICATE_db41 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1912_l1904_l1907_l1896_DUPLICATE_db41_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1907_c11_f74f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_9571 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_9571_return_output := result.is_stack_operation_16bit;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1904_l1920_l1907_l1896_DUPLICATE_0223 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1904_l1920_l1907_l1896_DUPLICATE_0223_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1920_c11_0923] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_left;
     BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_return_output := BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_398f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_398f_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1912_l1904_l1896_DUPLICATE_abe2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1912_l1904_l1896_DUPLICATE_abe2_return_output := result.is_sp_shift;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1904_l1907_l1896_DUPLICATE_68d6 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1904_l1907_l1896_DUPLICATE_68d6_return_output := result.sp_relative_shift;

     -- BIN_OP_DIV[uxn_opcodes_h_l1914_c26_c14d] LATENCY=0
     -- Inputs
     BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_left <= VAR_BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_left;
     BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_right <= VAR_BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_right;
     -- Outputs
     VAR_BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_return_output := BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1912_l1907_DUPLICATE_a08c LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1912_l1907_DUPLICATE_a08c_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_MUX_uxn_opcodes_h_l1914_c11_ba09_iffalse := VAR_BIN_OP_DIV_uxn_opcodes_h_l1914_c26_c14d_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1896_c2_257d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1896_c2_257d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1896_c6_819b_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1904_c11_d436_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1907_c11_f74f_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c11_e71f_return_output;
     VAR_MUX_uxn_opcodes_h_l1914_c11_ba09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1914_c11_9bf3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1920_c11_0923_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1904_l1907_l1896_DUPLICATE_68d6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1904_l1907_l1896_DUPLICATE_68d6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1904_l1907_l1896_DUPLICATE_68d6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1912_l1904_l1907_l1896_DUPLICATE_db41_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1912_l1904_l1907_l1896_DUPLICATE_db41_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1912_l1904_l1907_l1896_DUPLICATE_db41_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1912_l1904_l1907_l1896_DUPLICATE_db41_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_398f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_398f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_398f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_398f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1912_l1904_l1896_DUPLICATE_abe2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1912_l1904_l1896_DUPLICATE_abe2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1912_l1904_l1896_DUPLICATE_abe2_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_9571_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_9571_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_9571_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1912_l1904_l1920_l1907_DUPLICATE_9571_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1904_l1920_l1907_l1896_DUPLICATE_0223_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1904_l1920_l1907_l1896_DUPLICATE_0223_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1904_l1920_l1907_l1896_DUPLICATE_0223_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1904_l1920_l1907_l1896_DUPLICATE_0223_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1912_l1907_DUPLICATE_a08c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1912_l1907_DUPLICATE_a08c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_a0a9_return_output;
     -- t16_MUX[uxn_opcodes_h_l1907_c7_71a7] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond <= VAR_t16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond;
     t16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue;
     t16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output := t16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1920_c7_8e01] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output;

     -- n16_MUX[uxn_opcodes_h_l1912_c7_bb1d] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond <= VAR_n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond;
     n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue;
     n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output := n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1920_c7_8e01] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1912_c7_bb1d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1907_c7_71a7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;

     -- MUX[uxn_opcodes_h_l1914_c11_ba09] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1914_c11_ba09_cond <= VAR_MUX_uxn_opcodes_h_l1914_c11_ba09_cond;
     MUX_uxn_opcodes_h_l1914_c11_ba09_iftrue <= VAR_MUX_uxn_opcodes_h_l1914_c11_ba09_iftrue;
     MUX_uxn_opcodes_h_l1914_c11_ba09_iffalse <= VAR_MUX_uxn_opcodes_h_l1914_c11_ba09_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1914_c11_ba09_return_output := MUX_uxn_opcodes_h_l1914_c11_ba09_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1920_c7_8e01] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1912_c7_bb1d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;

     -- Submodule level 2
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue := VAR_MUX_uxn_opcodes_h_l1914_c11_ba09_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue := VAR_MUX_uxn_opcodes_h_l1914_c11_ba09_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1920_c7_8e01_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;
     -- t16_MUX[uxn_opcodes_h_l1904_c7_e7dd] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond <= VAR_t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond;
     t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue;
     t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output := t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1912_c7_bb1d] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1912_c7_bb1d] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond;
     tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output := tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1904_c7_e7dd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1912_c7_bb1d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1912_c7_bb1d] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output := result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1912_c7_bb1d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;

     -- n16_MUX[uxn_opcodes_h_l1907_c7_71a7] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond <= VAR_n16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond;
     n16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue;
     n16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output := n16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1907_c7_71a7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1907_c7_71a7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1912_c7_bb1d_return_output;
     -- n16_MUX[uxn_opcodes_h_l1904_c7_e7dd] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond <= VAR_n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond;
     n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue;
     n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output := n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1907_c7_71a7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;

     -- t16_MUX[uxn_opcodes_h_l1896_c2_257d] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1896_c2_257d_cond <= VAR_t16_MUX_uxn_opcodes_h_l1896_c2_257d_cond;
     t16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue;
     t16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output := t16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1907_c7_71a7] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_cond;
     tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output := tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1907_c7_71a7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1904_c7_e7dd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1896_c2_257d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1907_c7_71a7] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1904_c7_e7dd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1907_c7_71a7] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output := result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1907_c7_71a7_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1904_c7_e7dd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1896_c2_257d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1904_c7_e7dd] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output := result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1904_c7_e7dd] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;

     -- n16_MUX[uxn_opcodes_h_l1896_c2_257d] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1896_c2_257d_cond <= VAR_n16_MUX_uxn_opcodes_h_l1896_c2_257d_cond;
     n16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue;
     n16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output := n16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1904_c7_e7dd] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond;
     tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output := tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1896_c2_257d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1904_c7_e7dd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1904_c7_e7dd_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l1896_c2_257d] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_cond;
     tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output := tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1896_c2_257d] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_return_output := result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1896_c2_257d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1896_c2_257d] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1896_c2_257d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_return_output;

     -- Submodule level 6
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l1896_c2_257d_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1926_l1892_DUPLICATE_8d40 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1926_l1892_DUPLICATE_8d40_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1896_c2_257d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1896_c2_257d_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1926_l1892_DUPLICATE_8d40_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1926_l1892_DUPLICATE_8d40_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
