-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity nip2_0CLK_9a874500 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_9a874500;
architecture arch of nip2_0CLK_9a874500 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2053_c6_6d13]
signal BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2053_c1_7adc]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2053_c2_9f7a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2053_c2_9f7a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2053_c2_9f7a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2053_c2_9f7a]
signal result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2053_c2_9f7a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2053_c2_9f7a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2053_c2_9f7a]
signal t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l2054_c3_3492[uxn_opcodes_h_l2054_c3_3492]
signal printf_uxn_opcodes_h_l2054_c3_3492_uxn_opcodes_h_l2054_c3_3492_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2058_c11_f327]
signal BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2058_c7_fe78]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2058_c7_fe78]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2058_c7_fe78]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2058_c7_fe78]
signal result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2058_c7_fe78]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2058_c7_fe78]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2058_c7_fe78]
signal t16_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2061_c11_3481]
signal BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2061_c7_5bfd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2061_c7_5bfd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2061_c7_5bfd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2061_c7_5bfd]
signal result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2061_c7_5bfd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2061_c7_5bfd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2061_c7_5bfd]
signal t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2063_c3_2463]
signal CONST_SL_8_uxn_opcodes_h_l2063_c3_2463_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2063_c3_2463_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2065_c11_4cae]
signal BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2065_c7_13f5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2065_c7_13f5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2065_c7_13f5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2065_c7_13f5]
signal result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2065_c7_13f5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2065_c7_13f5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2065_c7_13f5]
signal t16_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2066_c3_e5c6]
signal BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2068_c30_9802]
signal sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2073_c11_7322]
signal BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2073_c7_9cd8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2073_c7_9cd8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2073_c7_9cd8]
signal result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2073_c7_9cd8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2073_c7_9cd8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output : unsigned(0 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l2076_c31_d2f7]
signal CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2078_c11_5167]
signal BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2078_c7_f5a7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2078_c7_f5a7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_c551( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13
BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_left,
BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_right,
BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a
result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a
result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a
result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a
result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output);

-- t16_MUX_uxn_opcodes_h_l2053_c2_9f7a
t16_MUX_uxn_opcodes_h_l2053_c2_9f7a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond,
t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue,
t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse,
t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output);

-- printf_uxn_opcodes_h_l2054_c3_3492_uxn_opcodes_h_l2054_c3_3492
printf_uxn_opcodes_h_l2054_c3_3492_uxn_opcodes_h_l2054_c3_3492 : entity work.printf_uxn_opcodes_h_l2054_c3_3492_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2054_c3_3492_uxn_opcodes_h_l2054_c3_3492_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327
BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_left,
BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_right,
BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78
result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78
result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78
result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_cond,
result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78
result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78
result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output);

-- t16_MUX_uxn_opcodes_h_l2058_c7_fe78
t16_MUX_uxn_opcodes_h_l2058_c7_fe78 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2058_c7_fe78_cond,
t16_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue,
t16_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse,
t16_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481
BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_left,
BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_right,
BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd
result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd
result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd
result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond,
result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd
result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd
result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output);

-- t16_MUX_uxn_opcodes_h_l2061_c7_5bfd
t16_MUX_uxn_opcodes_h_l2061_c7_5bfd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond,
t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue,
t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse,
t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2063_c3_2463
CONST_SL_8_uxn_opcodes_h_l2063_c3_2463 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2063_c3_2463_x,
CONST_SL_8_uxn_opcodes_h_l2063_c3_2463_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae
BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_left,
BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_right,
BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5
result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5
result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5
result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_cond,
result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5
result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5
result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output);

-- t16_MUX_uxn_opcodes_h_l2065_c7_13f5
t16_MUX_uxn_opcodes_h_l2065_c7_13f5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2065_c7_13f5_cond,
t16_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue,
t16_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse,
t16_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6
BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_left,
BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_right,
BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2068_c30_9802
sp_relative_shift_uxn_opcodes_h_l2068_c30_9802 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_ins,
sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_x,
sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_y,
sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322
BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_left,
BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_right,
BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8
result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8
result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8
result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8
result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output);

-- CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7
CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7_x,
CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167
BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_left,
BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_right,
BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7
result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output,
 t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output,
 t16_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output,
 t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output,
 CONST_SL_8_uxn_opcodes_h_l2063_c3_2463_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output,
 t16_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_return_output,
 sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output,
 CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2055_c3_505d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2054_c3_3492_uxn_opcodes_h_l2054_c3_3492_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2059_c3_981e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2058_c7_fe78_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2063_c3_2463_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2063_c3_2463_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2070_c3_8da1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2065_c7_13f5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_return_output : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2071_c21_2d97_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2075_c3_a9f7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2076_c21_0f43_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2058_l2053_l2078_l2073_DUPLICATE_a0fc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2053_l2065_l2058_l2061_DUPLICATE_03d1_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_6e92_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_b30b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2065_l2061_l2058_l2078_l2073_DUPLICATE_b1b6_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2062_l2066_DUPLICATE_197d_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2073_l2061_DUPLICATE_2f2a_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2083_l2049_DUPLICATE_f469_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2055_c3_505d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2055_c3_505d;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2075_c3_a9f7 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2075_c3_a9f7;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2070_c3_8da1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2070_c3_8da1;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2059_c3_981e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2059_c3_981e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_iffalse := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_left := t16;
     VAR_CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7_x := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l2078_c11_5167] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_left;
     BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_return_output := BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2053_l2065_l2058_l2061_DUPLICATE_03d1 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2053_l2065_l2058_l2061_DUPLICATE_03d1_return_output := result.sp_relative_shift;

     -- CONST_SR_8[uxn_opcodes_h_l2076_c31_d2f7] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7_x <= VAR_CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7_return_output := CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2058_l2053_l2078_l2073_DUPLICATE_a0fc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2058_l2053_l2078_l2073_DUPLICATE_a0fc_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2061_c11_3481] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_left;
     BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_return_output := BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2073_l2061_DUPLICATE_2f2a LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2073_l2061_DUPLICATE_2f2a_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l2068_c30_9802] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_ins;
     sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_x;
     sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_return_output := sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2065_c11_4cae] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_left;
     BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_return_output := BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2062_l2066_DUPLICATE_197d LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2062_l2066_DUPLICATE_197d_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l2058_c11_f327] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_left;
     BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_return_output := BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_b30b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_b30b_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2065_l2061_l2058_l2078_l2073_DUPLICATE_b1b6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2065_l2061_l2058_l2078_l2073_DUPLICATE_b1b6_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2073_c11_7322] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_left;
     BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_return_output := BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_6e92 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_6e92_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2053_c6_6d13] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_left;
     BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output := BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2053_c6_6d13_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2058_c7_fe78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2058_c11_f327_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c11_3481_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2065_c7_13f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2065_c11_4cae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_7322_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_5167_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2062_l2066_DUPLICATE_197d_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2063_c3_2463_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2062_l2066_DUPLICATE_197d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2053_l2065_l2058_l2061_DUPLICATE_03d1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2053_l2065_l2058_l2061_DUPLICATE_03d1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2053_l2065_l2058_l2061_DUPLICATE_03d1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2053_l2065_l2058_l2061_DUPLICATE_03d1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2065_l2061_l2058_l2078_l2073_DUPLICATE_b1b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2065_l2061_l2058_l2078_l2073_DUPLICATE_b1b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2065_l2061_l2058_l2078_l2073_DUPLICATE_b1b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2065_l2061_l2058_l2078_l2073_DUPLICATE_b1b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2065_l2061_l2058_l2078_l2073_DUPLICATE_b1b6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_b30b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_b30b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_b30b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_b30b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2058_l2053_l2078_l2073_DUPLICATE_a0fc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2058_l2053_l2078_l2073_DUPLICATE_a0fc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2058_l2053_l2078_l2073_DUPLICATE_a0fc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2058_l2053_l2078_l2073_DUPLICATE_a0fc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2058_l2053_l2078_l2073_DUPLICATE_a0fc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2073_l2061_DUPLICATE_2f2a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2073_l2061_DUPLICATE_2f2a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_6e92_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_6e92_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_6e92_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2053_l2058_l2073_l2061_DUPLICATE_6e92_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2068_c30_9802_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2073_c7_9cd8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2065_c7_13f5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2053_c1_7adc] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2078_c7_f5a7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2078_c7_f5a7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2073_c7_9cd8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2066_c3_e5c6] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_left;
     BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_return_output := BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2076_c21_0f43] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2076_c21_0f43_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l2076_c31_d2f7_return_output);

     -- CONST_SL_8[uxn_opcodes_h_l2063_c3_2463] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2063_c3_2463_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2063_c3_2463_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2063_c3_2463_return_output := CONST_SL_8_uxn_opcodes_h_l2063_c3_2463_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2076_c21_0f43_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2063_c3_2463_return_output;
     VAR_printf_uxn_opcodes_h_l2054_c3_3492_uxn_opcodes_h_l2054_c3_3492_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2053_c1_7adc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c7_f5a7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2065_c7_13f5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2073_c7_9cd8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2061_c7_5bfd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2073_c7_9cd8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output;

     -- printf_uxn_opcodes_h_l2054_c3_3492[uxn_opcodes_h_l2054_c3_3492] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2054_c3_3492_uxn_opcodes_h_l2054_c3_3492_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2054_c3_3492_uxn_opcodes_h_l2054_c3_3492_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2065_c7_13f5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;

     -- t16_MUX[uxn_opcodes_h_l2065_c7_13f5] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2065_c7_13f5_cond <= VAR_t16_MUX_uxn_opcodes_h_l2065_c7_13f5_cond;
     t16_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue;
     t16_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output := t16_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2071_c21_2d97] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2071_c21_2d97_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_BIN_OP_OR_uxn_opcodes_h_l2066_c3_e5c6_return_output);

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2073_c7_9cd8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2071_c21_2d97_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9cd8_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2065_c7_13f5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output := result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2058_c7_fe78] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2061_c7_5bfd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;

     -- t16_MUX[uxn_opcodes_h_l2061_c7_5bfd] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond <= VAR_t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond;
     t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue;
     t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output := t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2065_c7_13f5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2065_c7_13f5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2061_c7_5bfd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2065_c7_13f5_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2058_c7_fe78] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2061_c7_5bfd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output := result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2061_c7_5bfd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;

     -- t16_MUX[uxn_opcodes_h_l2058_c7_fe78] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2058_c7_fe78_cond <= VAR_t16_MUX_uxn_opcodes_h_l2058_c7_fe78_cond;
     t16_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue;
     t16_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output := t16_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2053_c2_9f7a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2061_c7_5bfd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2058_c7_fe78] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c7_5bfd_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2058_c7_fe78] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2053_c2_9f7a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2053_c2_9f7a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2058_c7_fe78] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;

     -- t16_MUX[uxn_opcodes_h_l2053_c2_9f7a] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond <= VAR_t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond;
     t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue;
     t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output := t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2058_c7_fe78] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output := result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2058_c7_fe78_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2053_c2_9f7a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2053_c2_9f7a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2053_c2_9f7a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2083_l2049_DUPLICATE_f469 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2083_l2049_DUPLICATE_f469_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c551(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2053_c2_9f7a_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2083_l2049_DUPLICATE_f469_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2083_l2049_DUPLICATE_f469_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
