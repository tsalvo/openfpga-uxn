-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 48
entity ldr_0CLK_f74745d5 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr_0CLK_f74745d5;
architecture arch of ldr_0CLK_f74745d5 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1599_c6_93ea]
signal BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1599_c2_4495]
signal t8_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1599_c2_4495]
signal tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1599_c2_4495]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1599_c2_4495]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1599_c2_4495]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1599_c2_4495]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1599_c2_4495]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1599_c2_4495]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1599_c2_4495]
signal result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1599_c2_4495]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1599_c2_4495]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1599_c2_4495]
signal result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1612_c11_d34f]
signal BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1612_c7_4b8f]
signal t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1612_c7_4b8f]
signal tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1612_c7_4b8f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : signed(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1612_c7_4b8f]
signal result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1612_c7_4b8f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1612_c7_4b8f]
signal result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1612_c7_4b8f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1612_c7_4b8f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1615_c11_fdfc]
signal BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1615_c7_aa7f]
signal t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1615_c7_aa7f]
signal tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1615_c7_aa7f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : signed(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1615_c7_aa7f]
signal result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1615_c7_aa7f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1615_c7_aa7f]
signal result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1615_c7_aa7f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1615_c7_aa7f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1617_c30_00e8]
signal sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1618_c22_ad01]
signal BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1620_c11_b15c]
signal BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1620_c7_1a45]
signal tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1620_c7_1a45]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1620_c7_1a45]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1620_c7_1a45]
signal result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1620_c7_1a45]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1620_c7_1a45]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1623_c11_3b7a]
signal BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1623_c7_9b3c]
signal tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1623_c7_9b3c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1623_c7_9b3c]
signal result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1623_c7_9b3c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1623_c7_9b3c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_d736( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.u16_value := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_vram_write := ref_toks_9;
      base.u8_value := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea
BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_left,
BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_right,
BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output);

-- t8_MUX_uxn_opcodes_h_l1599_c2_4495
t8_MUX_uxn_opcodes_h_l1599_c2_4495 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1599_c2_4495_cond,
t8_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue,
t8_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse,
t8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1599_c2_4495
tmp8_MUX_uxn_opcodes_h_l1599_c2_4495 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_cond,
tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue,
tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse,
tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495
result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495
result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495
result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495
result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495
result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_cond,
result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495
result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495
result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495
result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_cond,
result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f
BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_left,
BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_right,
BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output);

-- t8_MUX_uxn_opcodes_h_l1612_c7_4b8f
t8_MUX_uxn_opcodes_h_l1612_c7_4b8f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond,
t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue,
t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse,
t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f
tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond,
tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue,
tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse,
tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f
result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond,
result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f
result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f
result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f
result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc
BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_left,
BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_right,
BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output);

-- t8_MUX_uxn_opcodes_h_l1615_c7_aa7f
t8_MUX_uxn_opcodes_h_l1615_c7_aa7f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond,
t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue,
t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse,
t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f
tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond,
tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue,
tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse,
tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f
result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond,
result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f
result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f
result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8
sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_ins,
sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_x,
sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_y,
sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01
BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_left,
BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_right,
BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c
BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_left,
BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_right,
BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45
tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_cond,
tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue,
tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse,
tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45
result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45
result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45
result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_cond,
result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45
result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a
BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_left,
BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_right,
BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c
tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond,
tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue,
tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse,
tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c
result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c
result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c
result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output,
 t8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
 tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output,
 t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output,
 tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output,
 t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output,
 tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output,
 sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_return_output,
 tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_return_output,
 tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1604_c3_9c58 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1609_c3_59a1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1613_c3_7738 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1618_c3_7dd7 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1618_c27_fd65_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1621_c3_6b09 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1626_c3_ac46 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1615_l1599_l1612_DUPLICATE_444d_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1620_l1615_l1612_l1599_l1623_DUPLICATE_176c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1620_l1612_DUPLICATE_4c6a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_a75b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_32ea_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1615_l1620_l1623_DUPLICATE_76d2_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d736_uxn_opcodes_h_l1595_l1631_DUPLICATE_221c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1626_c3_ac46 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1626_c3_ac46;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1604_c3_9c58 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1604_c3_9c58;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_right := to_unsigned(2, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1613_c3_7738 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1613_c3_7738;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1609_c3_59a1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1609_c3_59a1;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1621_c3_6b09 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1621_c3_6b09;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1599_c6_93ea] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_left;
     BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output := BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1620_c11_b15c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1620_l1615_l1612_l1599_l1623_DUPLICATE_176c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1620_l1615_l1612_l1599_l1623_DUPLICATE_176c_return_output := result.u8_value;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1615_l1599_l1612_DUPLICATE_444d LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1615_l1599_l1612_DUPLICATE_444d_return_output := result.u16_value;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1599_c2_4495_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_a75b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_a75b_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1620_l1612_DUPLICATE_4c6a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1620_l1612_DUPLICATE_4c6a_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1623_c11_3b7a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1599_c2_4495_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_32ea LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_32ea_return_output := result.is_opc_done;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1599_c2_4495_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l1617_c30_00e8] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_ins;
     sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_x;
     sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_return_output := sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1612_c11_d34f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1618_c27_fd65] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1618_c27_fd65_return_output := CAST_TO_int8_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1615_c11_fdfc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_left;
     BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output := BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1599_c2_4495_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1615_l1620_l1623_DUPLICATE_76d2 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1615_l1620_l1623_DUPLICATE_76d2_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1599_c2_4495_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1599_c6_93ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_d34f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_fdfc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1620_c11_b15c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_3b7a_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1618_c27_fd65_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1620_l1612_DUPLICATE_4c6a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1620_l1612_DUPLICATE_4c6a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1615_l1599_l1612_DUPLICATE_444d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1615_l1599_l1612_DUPLICATE_444d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1615_l1599_l1612_DUPLICATE_444d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_32ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_32ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_32ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_32ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_a75b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_a75b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_a75b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1615_l1620_l1612_l1623_DUPLICATE_a75b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1615_l1620_l1623_DUPLICATE_76d2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1615_l1620_l1623_DUPLICATE_76d2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1615_l1620_l1623_DUPLICATE_76d2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1620_l1615_l1612_l1599_l1623_DUPLICATE_176c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1620_l1615_l1612_l1599_l1623_DUPLICATE_176c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1620_l1615_l1612_l1599_l1623_DUPLICATE_176c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1620_l1615_l1612_l1599_l1623_DUPLICATE_176c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1620_l1615_l1612_l1599_l1623_DUPLICATE_176c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1599_c2_4495_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1599_c2_4495_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1599_c2_4495_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1599_c2_4495_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1617_c30_00e8_return_output;
     -- BIN_OP_PLUS[uxn_opcodes_h_l1618_c22_ad01] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1623_c7_9b3c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1615_c7_aa7f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond;
     t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue;
     t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output := t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1623_c7_9b3c] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond;
     tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output := tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1623_c7_9b3c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1623_c7_9b3c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1620_c7_1a45] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1623_c7_9b3c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1618_c3_7dd7 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1618_c22_ad01_return_output)),16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1623_c7_9b3c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1618_c3_7dd7;
     -- result_u8_value_MUX[uxn_opcodes_h_l1620_c7_1a45] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output := result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1615_c7_aa7f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1620_c7_1a45] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_cond;
     tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output := tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1620_c7_1a45] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output;

     -- t8_MUX[uxn_opcodes_h_l1612_c7_4b8f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond;
     t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue;
     t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output := t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1620_c7_1a45] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1620_c7_1a45] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1615_c7_aa7f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output := result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1620_c7_1a45_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1615_c7_aa7f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1612_c7_4b8f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output := result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1612_c7_4b8f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1615_c7_aa7f] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond;
     tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output := tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1615_c7_aa7f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1599_c2_4495_cond <= VAR_t8_MUX_uxn_opcodes_h_l1599_c2_4495_cond;
     t8_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue;
     t8_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output := t8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1615_c7_aa7f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1615_c7_aa7f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1615_c7_aa7f_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output := result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1612_c7_4b8f] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond;
     tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output := tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1612_c7_4b8f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1612_c7_4b8f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1612_c7_4b8f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1612_c7_4b8f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1612_c7_4b8f_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output := result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1599_c2_4495] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_cond;
     tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output := tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;

     -- Submodule level 6
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1599_c2_4495_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_d736_uxn_opcodes_h_l1595_l1631_DUPLICATE_221c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d736_uxn_opcodes_h_l1595_l1631_DUPLICATE_221c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_d736(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1599_c2_4495_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1599_c2_4495_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d736_uxn_opcodes_h_l1595_l1631_DUPLICATE_221c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d736_uxn_opcodes_h_l1595_l1631_DUPLICATE_221c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
