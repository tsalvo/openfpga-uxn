-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 46
entity jsr_0CLK_fedec265 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr_0CLK_fedec265;
architecture arch of jsr_0CLK_fedec265 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l749_c6_06d9]
signal BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l749_c2_c884]
signal t8_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l749_c2_c884]
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l749_c2_c884]
signal result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l749_c2_c884]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l749_c2_c884]
signal result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l749_c2_c884]
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l749_c2_c884]
signal result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l749_c2_c884]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l749_c2_c884]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l749_c2_c884]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l749_c2_c884]
signal result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l762_c11_1421]
signal BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l762_c7_af4b]
signal t8_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l762_c7_af4b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l762_c7_af4b]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l762_c7_af4b]
signal result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l762_c7_af4b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l762_c7_af4b]
signal result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l762_c7_af4b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l762_c7_af4b]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l762_c7_af4b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l764_c30_7693]
signal sp_relative_shift_uxn_opcodes_h_l764_c30_7693_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l764_c30_7693_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l764_c30_7693_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l764_c30_7693_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l766_c11_4af1]
signal BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l766_c7_af0e]
signal t8_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l766_c7_af0e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l766_c7_af0e]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l766_c7_af0e]
signal result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l766_c7_af0e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l766_c7_af0e]
signal result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l766_c7_af0e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l766_c7_af0e]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l766_c7_af0e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l774_c11_c709]
signal BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l774_c7_7fcb]
signal result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l774_c7_7fcb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l774_c7_7fcb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l774_c7_7fcb]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l774_c7_7fcb]
signal result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l774_c7_7fcb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output : unsigned(0 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l777_c31_4e4f]
signal CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l779_c22_33bf]
signal BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_return_output : signed(17 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_775a( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.u16_value := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;
      base.is_ram_write := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9
BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_left,
BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_right,
BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output);

-- t8_MUX_uxn_opcodes_h_l749_c2_c884
t8_MUX_uxn_opcodes_h_l749_c2_c884 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l749_c2_c884_cond,
t8_MUX_uxn_opcodes_h_l749_c2_c884_iftrue,
t8_MUX_uxn_opcodes_h_l749_c2_c884_iffalse,
t8_MUX_uxn_opcodes_h_l749_c2_c884_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884
result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884
result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884
result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_cond,
result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884
result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884
result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_cond,
result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884
result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421
BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_left,
BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_right,
BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output);

-- t8_MUX_uxn_opcodes_h_l762_c7_af4b
t8_MUX_uxn_opcodes_h_l762_c7_af4b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l762_c7_af4b_cond,
t8_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue,
t8_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse,
t8_MUX_uxn_opcodes_h_l762_c7_af4b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b
result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b
result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_cond,
result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b
result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b
result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_cond,
result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b
result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b
result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l764_c30_7693
sp_relative_shift_uxn_opcodes_h_l764_c30_7693 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l764_c30_7693_ins,
sp_relative_shift_uxn_opcodes_h_l764_c30_7693_x,
sp_relative_shift_uxn_opcodes_h_l764_c30_7693_y,
sp_relative_shift_uxn_opcodes_h_l764_c30_7693_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1
BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_left,
BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_right,
BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output);

-- t8_MUX_uxn_opcodes_h_l766_c7_af0e
t8_MUX_uxn_opcodes_h_l766_c7_af0e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l766_c7_af0e_cond,
t8_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue,
t8_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse,
t8_MUX_uxn_opcodes_h_l766_c7_af0e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e
result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e
result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_cond,
result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e
result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e
result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_cond,
result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e
result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e
result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709
BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_left,
BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_right,
BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb
result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_cond,
result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb
result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb
result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb
result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_cond,
result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb
result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output);

-- CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f
CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f_x,
CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf
BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_left,
BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_right,
BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output,
 t8_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output,
 t8_MUX_uxn_opcodes_h_l762_c7_af4b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_return_output,
 sp_relative_shift_uxn_opcodes_h_l764_c30_7693_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output,
 t8_MUX_uxn_opcodes_h_l766_c7_af0e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output,
 CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l754_c3_9f54 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l759_c3_ad18 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l763_c3_5cc6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l764_c30_7693_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l764_c30_7693_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l764_c30_7693_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l764_c30_7693_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l769_c3_951c : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l771_c3_8bb5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l772_c21_4f35_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l779_c3_69d3 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l776_c3_9280 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l774_c7_7fcb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l775_c3_b263 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l774_c7_7fcb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l777_c21_766d_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l779_c27_48d2_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_return_output : signed(17 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l749_l762_l774_DUPLICATE_f00b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l749_l766_l762_l774_DUPLICATE_f39d_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l766_l762_DUPLICATE_d2f3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l766_l762_DUPLICATE_1e4f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l766_l762_l774_DUPLICATE_76b7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l766_l762_l774_DUPLICATE_42b6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_775a_uxn_opcodes_h_l783_l745_DUPLICATE_ebc3_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l764_c30_7693_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l754_c3_9f54 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l754_c3_9f54;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l771_c3_8bb5 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l771_c3_8bb5;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l776_c3_9280 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l776_c3_9280;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l759_c3_ad18 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l759_c3_ad18;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l769_c3_951c := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l769_c3_951c;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l775_c3_b263 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l775_c3_b263;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_right := to_unsigned(2, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l763_c3_5cc6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l763_c3_5cc6;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l764_c30_7693_y := resize(to_signed(-1, 2), 4);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l764_c30_7693_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f_x := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l749_c2_c884_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l766_l762_l774_DUPLICATE_76b7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l766_l762_l774_DUPLICATE_76b7_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l766_c11_4af1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_left;
     BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output := BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l749_c2_c884] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l749_c2_c884_return_output := result.is_ram_write;

     -- CONST_SR_8[uxn_opcodes_h_l777_c31_4e4f] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f_x <= VAR_CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f_return_output := CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l749_c6_06d9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_left;
     BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output := BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l749_l762_l774_DUPLICATE_f00b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l749_l762_l774_DUPLICATE_f00b_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l766_l762_DUPLICATE_d2f3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l766_l762_DUPLICATE_d2f3_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l749_l766_l762_l774_DUPLICATE_f39d LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l749_l766_l762_l774_DUPLICATE_f39d_return_output := result.u16_value;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l749_c2_c884] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l749_c2_c884_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l766_l762_DUPLICATE_1e4f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l766_l762_DUPLICATE_1e4f_return_output := result.is_stack_index_flipped;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l772_c21_4f35] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l772_c21_4f35_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_pc);

     -- sp_relative_shift[uxn_opcodes_h_l764_c30_7693] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l764_c30_7693_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l764_c30_7693_ins;
     sp_relative_shift_uxn_opcodes_h_l764_c30_7693_x <= VAR_sp_relative_shift_uxn_opcodes_h_l764_c30_7693_x;
     sp_relative_shift_uxn_opcodes_h_l764_c30_7693_y <= VAR_sp_relative_shift_uxn_opcodes_h_l764_c30_7693_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l764_c30_7693_return_output := sp_relative_shift_uxn_opcodes_h_l764_c30_7693_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l774_c7_7fcb] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l774_c7_7fcb_return_output := result.stack_address_sp_offset;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l774_c7_7fcb] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l774_c7_7fcb_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l762_c11_1421] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_left;
     BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output := BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l766_l762_l774_DUPLICATE_42b6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l766_l762_l774_DUPLICATE_42b6_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l774_c11_c709] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_left;
     BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_return_output := BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l779_c27_48d2] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l779_c27_48d2_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l749_c2_c884_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c6_06d9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l762_c7_af4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l762_c11_1421_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l766_c7_af0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l766_c11_4af1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l774_c11_c709_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l779_c27_48d2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l772_c21_4f35_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l749_l766_l762_l774_DUPLICATE_f39d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l749_l766_l762_l774_DUPLICATE_f39d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l749_l766_l762_l774_DUPLICATE_f39d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l749_l766_l762_l774_DUPLICATE_f39d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l766_l762_l774_DUPLICATE_76b7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l766_l762_l774_DUPLICATE_76b7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l766_l762_l774_DUPLICATE_76b7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l766_l762_l774_DUPLICATE_42b6_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l766_l762_l774_DUPLICATE_42b6_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l766_l762_l774_DUPLICATE_42b6_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l766_l762_DUPLICATE_1e4f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l766_l762_DUPLICATE_1e4f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l766_l762_DUPLICATE_d2f3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l766_l762_DUPLICATE_d2f3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l749_l762_l774_DUPLICATE_f00b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l749_l762_l774_DUPLICATE_f00b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l749_l762_l774_DUPLICATE_f00b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l749_c2_c884_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l749_c2_c884_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l774_c7_7fcb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l774_c7_7fcb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l764_c30_7693_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l774_c7_7fcb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l774_c7_7fcb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l774_c7_7fcb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l749_c2_c884] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l766_c7_af0e] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l766_c7_af0e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;

     -- t8_MUX[uxn_opcodes_h_l766_c7_af0e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l766_c7_af0e_cond <= VAR_t8_MUX_uxn_opcodes_h_l766_c7_af0e_cond;
     t8_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue;
     t8_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l766_c7_af0e_return_output := t8_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l749_c2_c884] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l779_c22_33bf] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_left;
     BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_return_output := BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l777_c21_766d] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l777_c21_766d_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l777_c31_4e4f_return_output);

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l774_c7_7fcb] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l779_c3_69d3 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l779_c22_33bf_return_output)),16);
     VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l777_c21_766d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue := VAR_result_u16_value_uxn_opcodes_h_l779_c3_69d3;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l762_c7_af4b] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l766_c7_af0e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l766_c7_af0e] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l774_c7_7fcb] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_cond;
     result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output := result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l766_c7_af0e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l766_c7_af0e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l762_c7_af4b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l774_c7_7fcb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output := result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output;

     -- t8_MUX[uxn_opcodes_h_l762_c7_af4b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l762_c7_af4b_cond <= VAR_t8_MUX_uxn_opcodes_h_l762_c7_af4b_cond;
     t8_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue;
     t8_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l762_c7_af4b_return_output := t8_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l774_c7_7fcb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l749_c2_c884_iffalse := VAR_t8_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l762_c7_af4b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l766_c7_af0e] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_cond;
     result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output := result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l762_c7_af4b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l766_c7_af0e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output := result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l762_c7_af4b] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;

     -- t8_MUX[uxn_opcodes_h_l749_c2_c884] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l749_c2_c884_cond <= VAR_t8_MUX_uxn_opcodes_h_l749_c2_c884_cond;
     t8_MUX_uxn_opcodes_h_l749_c2_c884_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l749_c2_c884_iftrue;
     t8_MUX_uxn_opcodes_h_l749_c2_c884_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l749_c2_c884_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l749_c2_c884_return_output := t8_MUX_uxn_opcodes_h_l749_c2_c884_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l749_c2_c884] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l762_c7_af4b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l749_c2_c884] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l766_c7_af0e_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l749_c2_c884_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l749_c2_c884] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l749_c2_c884] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l749_c2_c884] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l749_c2_c884] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l762_c7_af4b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output := result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l762_c7_af4b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output := result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;

     -- Submodule level 5
     VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l762_c7_af4b_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l749_c2_c884] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_cond;
     result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output := result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l749_c2_c884] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_cond;
     result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output := result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_775a_uxn_opcodes_h_l783_l745_DUPLICATE_ebc3 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_775a_uxn_opcodes_h_l783_l745_DUPLICATE_ebc3_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_775a(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c2_c884_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l749_c2_c884_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_775a_uxn_opcodes_h_l783_l745_DUPLICATE_ebc3_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_775a_uxn_opcodes_h_l783_l745_DUPLICATE_ebc3_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
