-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity ldz_0CLK_f74745d5 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_f74745d5;
architecture arch of ldz_0CLK_f74745d5 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1521_c6_ccbd]
signal BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1521_c2_0faa]
signal tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1521_c2_0faa]
signal t8_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1521_c2_0faa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1521_c2_0faa]
signal result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1521_c2_0faa]
signal result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1521_c2_0faa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1521_c2_0faa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1521_c2_0faa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1521_c2_0faa]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1526_c11_7ef5]
signal BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1526_c7_2f8e]
signal tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1526_c7_2f8e]
signal t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1526_c7_2f8e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1526_c7_2f8e]
signal result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1526_c7_2f8e]
signal result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1526_c7_2f8e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1526_c7_2f8e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1526_c7_2f8e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1526_c7_2f8e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1529_c11_a7ec]
signal BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1529_c7_184a]
signal tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1529_c7_184a]
signal t8_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1529_c7_184a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1529_c7_184a]
signal result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1529_c7_184a]
signal result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1529_c7_184a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1529_c7_184a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1529_c7_184a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1529_c7_184a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1532_c30_d857]
signal sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1535_c11_6161]
signal BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1535_c7_5ff5]
signal tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1535_c7_5ff5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1535_c7_5ff5]
signal result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1535_c7_5ff5]
signal result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1535_c7_5ff5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1535_c7_5ff5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1535_c7_5ff5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1539_c11_a1c7]
signal BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1539_c7_9265]
signal tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1539_c7_9265]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1539_c7_9265]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1539_c7_9265]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1539_c7_9265]
signal result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1545_c11_fdc0]
signal BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1545_c7_8e4a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1545_c7_8e4a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_sp_shift := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd
BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_left,
BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_right,
BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa
tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_cond,
tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue,
tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse,
tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output);

-- t8_MUX_uxn_opcodes_h_l1521_c2_0faa
t8_MUX_uxn_opcodes_h_l1521_c2_0faa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1521_c2_0faa_cond,
t8_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue,
t8_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse,
t8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa
result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_cond,
result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa
result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_cond,
result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa
result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa
result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa
result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa
result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5
BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_left,
BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_right,
BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e
tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond,
tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue,
tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse,
tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output);

-- t8_MUX_uxn_opcodes_h_l1526_c7_2f8e
t8_MUX_uxn_opcodes_h_l1526_c7_2f8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond,
t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue,
t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse,
t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e
result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e
result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond,
result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e
result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e
result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e
result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec
BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_left,
BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_right,
BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1529_c7_184a
tmp8_MUX_uxn_opcodes_h_l1529_c7_184a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_cond,
tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue,
tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse,
tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output);

-- t8_MUX_uxn_opcodes_h_l1529_c7_184a
t8_MUX_uxn_opcodes_h_l1529_c7_184a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1529_c7_184a_cond,
t8_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue,
t8_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse,
t8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a
result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a
result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_cond,
result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a
result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a
result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a
result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1532_c30_d857
sp_relative_shift_uxn_opcodes_h_l1532_c30_d857 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_ins,
sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_x,
sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_y,
sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161
BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_left,
BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_right,
BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5
tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond,
tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue,
tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse,
tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5
result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5
result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond,
result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5
result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5
result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5
result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7
BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_left,
BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_right,
BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1539_c7_9265
tmp8_MUX_uxn_opcodes_h_l1539_c7_9265 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_cond,
tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue,
tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse,
tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265
result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265
result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265
result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_cond,
result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0
BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_left,
BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_right,
BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a
result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a
result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output,
 tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
 t8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output,
 tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output,
 t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output,
 tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output,
 t8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output,
 sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_return_output,
 tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_return_output,
 tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1523_c3_360a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1527_c3_8eeb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1533_c22_49c9_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1537_c22_4c87_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1542_c3_da34 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1539_DUPLICATE_2c91_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1521_l1535_l1526_DUPLICATE_8c82_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1545_DUPLICATE_49cf_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1529_l1521_l1526_DUPLICATE_70dc_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1521_l1535_l1526_DUPLICATE_2ee4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1545_l1539_DUPLICATE_02a7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1529_l1539_l1535_DUPLICATE_5496_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce_uxn_opcodes_h_l1517_l1550_DUPLICATE_3073_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1542_c3_da34 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1542_c3_da34;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1523_c3_360a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1523_c3_360a;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1527_c3_8eeb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1527_c3_8eeb;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse := tmp8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1545_l1539_DUPLICATE_02a7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1545_l1539_DUPLICATE_02a7_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1521_l1535_l1526_DUPLICATE_2ee4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1521_l1535_l1526_DUPLICATE_2ee4_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1529_l1539_l1535_DUPLICATE_5496 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1529_l1539_l1535_DUPLICATE_5496_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1521_c6_ccbd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_left;
     BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output := BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1529_l1521_l1526_DUPLICATE_70dc LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1529_l1521_l1526_DUPLICATE_70dc_return_output := result.sp_relative_shift;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1533_c22_49c9] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1533_c22_49c9_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1537_c22_4c87] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1537_c22_4c87_return_output := CAST_TO_uint16_t_uint8_t(
     t8);

     -- BIN_OP_EQ[uxn_opcodes_h_l1526_c11_7ef5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1539_c11_a1c7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_left;
     BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_return_output := BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1535_c11_6161] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_left;
     BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_return_output := BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1545_DUPLICATE_49cf LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1545_DUPLICATE_49cf_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1529_c11_a7ec] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_left;
     BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output := BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1532_c30_d857] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_ins;
     sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_x;
     sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_return_output := sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1545_c11_fdc0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1521_l1535_l1526_DUPLICATE_8c82 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1521_l1535_l1526_DUPLICATE_8c82_return_output := result.u16_value;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1539_DUPLICATE_2c91 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1539_DUPLICATE_2c91_return_output := result.u8_value;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1521_c2_0faa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1521_c6_ccbd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_7ef5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1529_c7_184a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a7ec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_6161_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1539_c11_a1c7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1545_c11_fdc0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1533_c22_49c9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1537_c22_4c87_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1529_l1521_l1526_DUPLICATE_70dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1529_l1521_l1526_DUPLICATE_70dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1529_l1521_l1526_DUPLICATE_70dc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1521_l1535_l1526_DUPLICATE_8c82_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1521_l1535_l1526_DUPLICATE_8c82_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1521_l1535_l1526_DUPLICATE_8c82_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1545_l1539_DUPLICATE_02a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1545_l1539_DUPLICATE_02a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1545_l1539_DUPLICATE_02a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1545_l1539_DUPLICATE_02a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1545_l1539_DUPLICATE_02a7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1521_l1535_l1526_DUPLICATE_2ee4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1521_l1535_l1526_DUPLICATE_2ee4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1521_l1535_l1526_DUPLICATE_2ee4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1545_DUPLICATE_49cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1545_DUPLICATE_49cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1545_DUPLICATE_49cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1545_DUPLICATE_49cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1545_DUPLICATE_49cf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1529_l1539_l1535_DUPLICATE_5496_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1529_l1539_l1535_DUPLICATE_5496_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1529_l1539_l1535_DUPLICATE_5496_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1539_DUPLICATE_2c91_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1539_DUPLICATE_2c91_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1539_DUPLICATE_2c91_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1539_DUPLICATE_2c91_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1535_l1529_l1526_l1521_l1539_DUPLICATE_2c91_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1532_c30_d857_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1545_c7_8e4a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1535_c7_5ff5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1539_c7_9265] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1539_c7_9265] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_cond;
     tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_return_output := tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1535_c7_5ff5] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output := result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;

     -- t8_MUX[uxn_opcodes_h_l1529_c7_184a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1529_c7_184a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1529_c7_184a_cond;
     t8_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue;
     t8_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output := t8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1529_c7_184a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1539_c7_9265] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_return_output := result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1545_c7_8e4a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1545_c7_8e4a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1539_c7_9265_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1539_c7_9265_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1539_c7_9265_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1529_c7_184a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1535_c7_5ff5] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond;
     tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output := tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1535_c7_5ff5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1529_c7_184a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output := result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1535_c7_5ff5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1539_c7_9265] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_return_output;

     -- t8_MUX[uxn_opcodes_h_l1526_c7_2f8e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond <= VAR_t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond;
     t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue;
     t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output := t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1539_c7_9265] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1526_c7_2f8e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1539_c7_9265_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1539_c7_9265_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1526_c7_2f8e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1535_c7_5ff5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1529_c7_184a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1535_c7_5ff5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1526_c7_2f8e] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output := result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1521_c2_0faa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output;

     -- t8_MUX[uxn_opcodes_h_l1521_c2_0faa] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1521_c2_0faa_cond <= VAR_t8_MUX_uxn_opcodes_h_l1521_c2_0faa_cond;
     t8_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue;
     t8_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output := t8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1529_c7_184a] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_cond;
     tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output := tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1529_c7_184a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1535_c7_5ff5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1526_c7_2f8e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1529_c7_184a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1526_c7_2f8e] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond;
     tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output := tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1521_c2_0faa] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output := result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1529_c7_184a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1521_c2_0faa] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1526_c7_2f8e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_184a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1521_c2_0faa] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output := result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1526_c7_2f8e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1521_c2_0faa] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_cond;
     tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output := tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1521_c2_0faa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1526_c7_2f8e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_2f8e_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1521_c2_0faa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1521_c2_0faa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce_uxn_opcodes_h_l1517_l1550_DUPLICATE_3073 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce_uxn_opcodes_h_l1517_l1550_DUPLICATE_3073_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1521_c2_0faa_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce_uxn_opcodes_h_l1517_l1550_DUPLICATE_3073_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b7ce_uxn_opcodes_h_l1517_l1550_DUPLICATE_3073_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
