-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 46
entity jsr_0CLK_fedec265 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr_0CLK_fedec265;
architecture arch of jsr_0CLK_fedec265 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l754_c6_9d57]
signal BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l754_c2_dc3c]
signal t8_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l754_c2_dc3c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l754_c2_dc3c]
signal result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l754_c2_dc3c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l754_c2_dc3c]
signal result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l754_c2_dc3c]
signal result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l754_c2_dc3c]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l754_c2_dc3c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l754_c2_dc3c]
signal result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l754_c2_dc3c]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l754_c2_dc3c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l767_c11_d9d0]
signal BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l767_c7_ecc3]
signal t8_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l767_c7_ecc3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l767_c7_ecc3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l767_c7_ecc3]
signal result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l767_c7_ecc3]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l767_c7_ecc3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l767_c7_ecc3]
signal result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l767_c7_ecc3]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l767_c7_ecc3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l769_c30_8a4c]
signal sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l771_c11_a85c]
signal BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l771_c7_4816]
signal t8_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l771_c7_4816]
signal result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l771_c7_4816]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l771_c7_4816]
signal result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l771_c7_4816]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l771_c7_4816]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l771_c7_4816]
signal result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l771_c7_4816]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l771_c7_4816]
signal result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l779_c11_f6ab]
signal BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l779_c7_343d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l779_c7_343d]
signal result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l779_c7_343d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l779_c7_343d]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l779_c7_343d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l779_c7_343d]
signal result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output : unsigned(7 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l782_c31_26ac]
signal CONST_SR_8_uxn_opcodes_h_l782_c31_26ac_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l782_c31_26ac_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l784_c22_ca52]
signal BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_return_output : signed(17 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.u16_value := ref_toks_8;
      base.is_pc_updated := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57
BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_left,
BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_right,
BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output);

-- t8_MUX_uxn_opcodes_h_l754_c2_dc3c
t8_MUX_uxn_opcodes_h_l754_c2_dc3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l754_c2_dc3c_cond,
t8_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue,
t8_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse,
t8_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c
result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c
result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c
result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c
result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_cond,
result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c
result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_cond,
result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c
result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0
BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_left,
BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_right,
BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output);

-- t8_MUX_uxn_opcodes_h_l767_c7_ecc3
t8_MUX_uxn_opcodes_h_l767_c7_ecc3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l767_c7_ecc3_cond,
t8_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue,
t8_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse,
t8_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3
result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3
result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3
result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_cond,
result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3
result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_cond,
result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3
result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3
result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output);

-- sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c
sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_ins,
sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_x,
sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_y,
sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c
BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_left,
BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_right,
BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output);

-- t8_MUX_uxn_opcodes_h_l771_c7_4816
t8_MUX_uxn_opcodes_h_l771_c7_4816 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l771_c7_4816_cond,
t8_MUX_uxn_opcodes_h_l771_c7_4816_iftrue,
t8_MUX_uxn_opcodes_h_l771_c7_4816_iffalse,
t8_MUX_uxn_opcodes_h_l771_c7_4816_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816
result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816
result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816
result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_cond,
result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816
result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_cond,
result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816
result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816
result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab
BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_left,
BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_right,
BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d
result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_cond,
result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d
result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d
result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d
result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d
result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_cond,
result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output);

-- CONST_SR_8_uxn_opcodes_h_l782_c31_26ac
CONST_SR_8_uxn_opcodes_h_l782_c31_26ac : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l782_c31_26ac_x,
CONST_SR_8_uxn_opcodes_h_l782_c31_26ac_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52
BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_left,
BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_right,
BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output,
 t8_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output,
 t8_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output,
 sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output,
 t8_MUX_uxn_opcodes_h_l771_c7_4816_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output,
 CONST_SR_8_uxn_opcodes_h_l782_c31_26ac_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l759_c3_f13c : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l764_c3_88d2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l768_c3_4189 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l774_c3_f8f7 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l776_c3_15d6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l777_c21_e6a2_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l781_c3_854d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l779_c7_343d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l784_c3_a421 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l780_c3_04d8 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l779_c7_343d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l782_c31_26ac_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l782_c31_26ac_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l782_c21_6b57_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l784_c27_9551_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_return_output : signed(17 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l754_l779_l767_DUPLICATE_e0e1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l771_l754_l779_l767_DUPLICATE_73ce_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l771_l767_DUPLICATE_444e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l771_l767_DUPLICATE_701e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l771_l779_l767_DUPLICATE_8218_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l771_l779_l767_DUPLICATE_9ca1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l788_l750_DUPLICATE_5e33_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l768_c3_4189 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l768_c3_4189;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l764_c3_88d2 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l764_c3_88d2;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l774_c3_f8f7 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l774_c3_f8f7;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l776_c3_15d6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l776_c3_15d6;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l781_c3_854d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l781_c3_854d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_right := to_unsigned(3, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l759_c3_f13c := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l759_c3_f13c;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l780_c3_04d8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l780_c3_04d8;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_CONST_SR_8_uxn_opcodes_h_l782_c31_26ac_x := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l771_c7_4816_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l771_c7_4816_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l769_c30_8a4c] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_ins;
     sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_x <= VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_x;
     sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_y <= VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_return_output := sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l771_l767_DUPLICATE_444e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l771_l767_DUPLICATE_444e_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l767_c11_d9d0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_left;
     BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output := BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l754_c2_dc3c] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l754_c2_dc3c_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l771_l767_DUPLICATE_701e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l771_l767_DUPLICATE_701e_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l771_l779_l767_DUPLICATE_8218 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l771_l779_l767_DUPLICATE_8218_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l754_c6_9d57] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_left;
     BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output := BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l754_l779_l767_DUPLICATE_e0e1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l754_l779_l767_DUPLICATE_e0e1_return_output := result.u8_value;

     -- CAST_TO_int8_t[uxn_opcodes_h_l784_c27_9551] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l784_c27_9551_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- CONST_SR_8[uxn_opcodes_h_l782_c31_26ac] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l782_c31_26ac_x <= VAR_CONST_SR_8_uxn_opcodes_h_l782_c31_26ac_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l782_c31_26ac_return_output := CONST_SR_8_uxn_opcodes_h_l782_c31_26ac_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l754_c2_dc3c] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l754_c2_dc3c_return_output := result.is_ram_write;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l777_c21_e6a2] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l777_c21_e6a2_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_pc);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l771_l779_l767_DUPLICATE_9ca1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l771_l779_l767_DUPLICATE_9ca1_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l771_l754_l779_l767_DUPLICATE_73ce LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l771_l754_l779_l767_DUPLICATE_73ce_return_output := result.u16_value;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l779_c7_343d] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l779_c7_343d_return_output := result.sp_relative_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l779_c7_343d] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l779_c7_343d_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l771_c11_a85c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_left;
     BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output := BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l779_c11_f6ab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_left;
     BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_return_output := BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l754_c2_dc3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9d57_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l767_c7_ecc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_d9d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l771_c7_4816_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_a85c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_f6ab_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l784_c27_9551_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l777_c21_e6a2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l771_l754_l779_l767_DUPLICATE_73ce_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l771_l754_l779_l767_DUPLICATE_73ce_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l771_l754_l779_l767_DUPLICATE_73ce_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l771_l754_l779_l767_DUPLICATE_73ce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l771_l779_l767_DUPLICATE_9ca1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l771_l779_l767_DUPLICATE_9ca1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l771_l779_l767_DUPLICATE_9ca1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l771_l779_l767_DUPLICATE_8218_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l771_l779_l767_DUPLICATE_8218_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l771_l779_l767_DUPLICATE_8218_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l771_l767_DUPLICATE_701e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l771_l767_DUPLICATE_701e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l771_l767_DUPLICATE_444e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l771_l767_DUPLICATE_444e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l754_l779_l767_DUPLICATE_e0e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l754_l779_l767_DUPLICATE_e0e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l754_l779_l767_DUPLICATE_e0e1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l754_c2_dc3c_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l754_c2_dc3c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l779_c7_343d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l779_c7_343d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_8a4c_return_output;
     -- t8_MUX[uxn_opcodes_h_l771_c7_4816] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l771_c7_4816_cond <= VAR_t8_MUX_uxn_opcodes_h_l771_c7_4816_cond;
     t8_MUX_uxn_opcodes_h_l771_c7_4816_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l771_c7_4816_iftrue;
     t8_MUX_uxn_opcodes_h_l771_c7_4816_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l771_c7_4816_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l771_c7_4816_return_output := t8_MUX_uxn_opcodes_h_l771_c7_4816_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l779_c7_343d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l784_c22_ca52] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_left;
     BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_return_output := BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l782_c21_6b57] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l782_c21_6b57_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l782_c31_26ac_return_output);

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l779_c7_343d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l771_c7_4816] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l754_c2_dc3c] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l779_c7_343d] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l771_c7_4816] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l754_c2_dc3c] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l779_c7_343d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l784_c3_a421 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_ca52_return_output)),16);
     VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l782_c21_6b57_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_343d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_343d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_4816_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_4816_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_343d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_343d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse := VAR_t8_MUX_uxn_opcodes_h_l771_c7_4816_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_iftrue := VAR_result_u16_value_uxn_opcodes_h_l784_c3_a421;
     -- result_u8_value_MUX[uxn_opcodes_h_l779_c7_343d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output := result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l771_c7_4816] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l771_c7_4816] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l771_c7_4816] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l767_c7_ecc3] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l779_c7_343d] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_cond;
     result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output := result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l771_c7_4816] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_return_output;

     -- t8_MUX[uxn_opcodes_h_l767_c7_ecc3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l767_c7_ecc3_cond <= VAR_t8_MUX_uxn_opcodes_h_l767_c7_ecc3_cond;
     t8_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue;
     t8_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output := t8_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l767_c7_ecc3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_4816_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_4816_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_4816_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_4816_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_343d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l767_c7_ecc3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l771_c7_4816] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_cond;
     result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output := result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l767_c7_ecc3] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l754_c2_dc3c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l767_c7_ecc3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;

     -- t8_MUX[uxn_opcodes_h_l754_c2_dc3c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l754_c2_dc3c_cond <= VAR_t8_MUX_uxn_opcodes_h_l754_c2_dc3c_cond;
     t8_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue;
     t8_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output := t8_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l754_c2_dc3c] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l771_c7_4816] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_cond;
     result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output := result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l767_c7_ecc3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_4816_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l754_c2_dc3c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l754_c2_dc3c] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l754_c2_dc3c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l767_c7_ecc3] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_cond;
     result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output := result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l767_c7_ecc3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output := result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l754_c2_dc3c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output;

     -- Submodule level 5
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_ecc3_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l754_c2_dc3c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output := result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l754_c2_dc3c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output := result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l788_l750_DUPLICATE_5e33 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l788_l750_DUPLICATE_5e33_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_dc3c_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l788_l750_DUPLICATE_5e33_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l788_l750_DUPLICATE_5e33_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
