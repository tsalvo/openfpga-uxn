-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 42
entity swp_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end swp_0CLK_64d180f1;
architecture arch of swp_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2508_c6_825e]
signal BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2508_c2_0684]
signal n8_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2508_c2_0684]
signal result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2508_c2_0684]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2508_c2_0684]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2508_c2_0684]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2508_c2_0684]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2508_c2_0684]
signal t8_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2515_c11_c3cd]
signal BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2515_c7_f90d]
signal n8_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2515_c7_f90d]
signal result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2515_c7_f90d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2515_c7_f90d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2515_c7_f90d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2515_c7_f90d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2515_c7_f90d]
signal t8_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2518_c11_699a]
signal BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2518_c7_09c2]
signal n8_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2518_c7_09c2]
signal result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2518_c7_09c2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2518_c7_09c2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2518_c7_09c2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2518_c7_09c2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2518_c7_09c2]
signal t8_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2521_c11_f4d8]
signal BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2521_c7_f6be]
signal n8_MUX_uxn_opcodes_h_l2521_c7_f6be_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2521_c7_f6be]
signal result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2521_c7_f6be]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2521_c7_f6be]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2521_c7_f6be]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2521_c7_f6be]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2524_c30_e2f3]
signal sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2529_c11_2fe2]
signal BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2529_c7_5cbd]
signal result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2529_c7_5cbd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2529_c7_5cbd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2529_c7_5cbd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2529_c7_5cbd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2534_c11_516d]
signal BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2534_c7_d51e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2534_c7_d51e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e
BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_left,
BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_right,
BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_return_output);

-- n8_MUX_uxn_opcodes_h_l2508_c2_0684
n8_MUX_uxn_opcodes_h_l2508_c2_0684 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2508_c2_0684_cond,
n8_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue,
n8_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse,
n8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684
result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_cond,
result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684
result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684
result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684
result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_return_output);

-- t8_MUX_uxn_opcodes_h_l2508_c2_0684
t8_MUX_uxn_opcodes_h_l2508_c2_0684 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2508_c2_0684_cond,
t8_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue,
t8_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse,
t8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd
BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_left,
BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_right,
BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_return_output);

-- n8_MUX_uxn_opcodes_h_l2515_c7_f90d
n8_MUX_uxn_opcodes_h_l2515_c7_f90d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2515_c7_f90d_cond,
n8_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue,
n8_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse,
n8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d
result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d
result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d
result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output);

-- t8_MUX_uxn_opcodes_h_l2515_c7_f90d
t8_MUX_uxn_opcodes_h_l2515_c7_f90d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2515_c7_f90d_cond,
t8_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue,
t8_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse,
t8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a
BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_left,
BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_right,
BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_return_output);

-- n8_MUX_uxn_opcodes_h_l2518_c7_09c2
n8_MUX_uxn_opcodes_h_l2518_c7_09c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2518_c7_09c2_cond,
n8_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue,
n8_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse,
n8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2
result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2
result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2
result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output);

-- t8_MUX_uxn_opcodes_h_l2518_c7_09c2
t8_MUX_uxn_opcodes_h_l2518_c7_09c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2518_c7_09c2_cond,
t8_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue,
t8_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse,
t8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8
BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_left,
BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_right,
BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_return_output);

-- n8_MUX_uxn_opcodes_h_l2521_c7_f6be
n8_MUX_uxn_opcodes_h_l2521_c7_f6be : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2521_c7_f6be_cond,
n8_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue,
n8_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse,
n8_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be
result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_cond,
result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be
result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be
result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be
result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3
sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_ins,
sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_x,
sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_y,
sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2
BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_left,
BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_right,
BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd
result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond,
result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd
result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd
result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd
result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d
BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_left,
BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_right,
BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e
result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e
result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_return_output,
 n8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_return_output,
 t8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_return_output,
 n8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output,
 t8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_return_output,
 n8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output,
 t8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_return_output,
 n8_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output,
 sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2512_c3_73dd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2508_c2_0684_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2516_c3_f09a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2515_c7_f90d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2518_c7_09c2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2521_c7_f6be_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2526_c3_f4f2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2531_c3_60cb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2530_c3_6413 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_bc11_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2508_l2534_l2529_l2518_l2515_DUPLICATE_7d6b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_8daf_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2534_l2529_l2521_l2518_l2515_DUPLICATE_2d10_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2529_l2518_DUPLICATE_63e3_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2539_l2504_DUPLICATE_99f5_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2530_c3_6413 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2530_c3_6413;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2512_c3_73dd := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2512_c3_73dd;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2531_c3_60cb := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2531_c3_60cb;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2526_c3_f4f2 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2526_c3_f4f2;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2516_c3_f09a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2516_c3_f09a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse := t8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2529_l2518_DUPLICATE_63e3 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2529_l2518_DUPLICATE_63e3_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2534_l2529_l2521_l2518_l2515_DUPLICATE_2d10 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2534_l2529_l2521_l2518_l2515_DUPLICATE_2d10_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2521_c11_f4d8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2518_c11_699a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2515_c11_c3cd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2534_c11_516d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_bc11 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_bc11_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_8daf LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_8daf_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l2524_c30_e2f3] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_ins;
     sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_x;
     sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_return_output := sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2508_l2534_l2529_l2518_l2515_DUPLICATE_7d6b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2508_l2534_l2529_l2518_l2515_DUPLICATE_7d6b_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2529_c11_2fe2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2508_c6_825e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2508_c2_0684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2508_c2_0684_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2508_c6_825e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2515_c7_f90d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2515_c7_f90d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2515_c11_c3cd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2518_c7_09c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2518_c7_09c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2518_c11_699a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2521_c7_f6be_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2521_c11_f4d8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2529_c11_2fe2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2534_c11_516d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_8daf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_8daf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_8daf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_8daf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2534_l2529_l2521_l2518_l2515_DUPLICATE_2d10_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2534_l2529_l2521_l2518_l2515_DUPLICATE_2d10_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2534_l2529_l2521_l2518_l2515_DUPLICATE_2d10_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2534_l2529_l2521_l2518_l2515_DUPLICATE_2d10_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2534_l2529_l2521_l2518_l2515_DUPLICATE_2d10_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2508_l2534_l2529_l2518_l2515_DUPLICATE_7d6b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2508_l2534_l2529_l2518_l2515_DUPLICATE_7d6b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2508_l2534_l2529_l2518_l2515_DUPLICATE_7d6b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2508_l2534_l2529_l2518_l2515_DUPLICATE_7d6b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2508_l2534_l2529_l2518_l2515_DUPLICATE_7d6b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2529_l2518_DUPLICATE_63e3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2529_l2518_DUPLICATE_63e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_bc11_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_bc11_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_bc11_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2508_l2515_l2529_l2518_DUPLICATE_bc11_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2524_c30_e2f3_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2529_c7_5cbd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2529_c7_5cbd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output;

     -- n8_MUX[uxn_opcodes_h_l2521_c7_f6be] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2521_c7_f6be_cond <= VAR_n8_MUX_uxn_opcodes_h_l2521_c7_f6be_cond;
     n8_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue;
     n8_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output := n8_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2534_c7_d51e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2534_c7_d51e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output;

     -- t8_MUX[uxn_opcodes_h_l2518_c7_09c2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2518_c7_09c2_cond <= VAR_t8_MUX_uxn_opcodes_h_l2518_c7_09c2_cond;
     t8_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue;
     t8_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output := t8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2529_c7_5cbd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output := result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2534_c7_d51e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2529_c7_5cbd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2521_c7_f6be] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2529_c7_5cbd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output;

     -- t8_MUX[uxn_opcodes_h_l2515_c7_f90d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2515_c7_f90d_cond <= VAR_t8_MUX_uxn_opcodes_h_l2515_c7_f90d_cond;
     t8_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue;
     t8_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output := t8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2521_c7_f6be] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output := result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2521_c7_f6be] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output;

     -- n8_MUX[uxn_opcodes_h_l2518_c7_09c2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2518_c7_09c2_cond <= VAR_n8_MUX_uxn_opcodes_h_l2518_c7_09c2_cond;
     n8_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue;
     n8_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output := n8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2529_c7_5cbd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;
     -- t8_MUX[uxn_opcodes_h_l2508_c2_0684] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2508_c2_0684_cond <= VAR_t8_MUX_uxn_opcodes_h_l2508_c2_0684_cond;
     t8_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue;
     t8_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output := t8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2518_c7_09c2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2521_c7_f6be] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2518_c7_09c2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2518_c7_09c2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;

     -- n8_MUX[uxn_opcodes_h_l2515_c7_f90d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2515_c7_f90d_cond <= VAR_n8_MUX_uxn_opcodes_h_l2515_c7_f90d_cond;
     n8_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue;
     n8_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output := n8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2521_c7_f6be] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2521_c7_f6be_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2518_c7_09c2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2515_c7_f90d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2515_c7_f90d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2515_c7_f90d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;

     -- n8_MUX[uxn_opcodes_h_l2508_c2_0684] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2508_c2_0684_cond <= VAR_n8_MUX_uxn_opcodes_h_l2508_c2_0684_cond;
     n8_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue;
     n8_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output := n8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2518_c7_09c2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2508_c2_0684_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2518_c7_09c2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2515_c7_f90d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2508_c2_0684] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2515_c7_f90d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2508_c2_0684] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2508_c2_0684] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_return_output := result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2515_c7_f90d_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2508_c2_0684] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2508_c2_0684] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2539_l2504_DUPLICATE_99f5 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2539_l2504_DUPLICATE_99f5_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2508_c2_0684_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2508_c2_0684_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2508_c2_0684_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2508_c2_0684_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2508_c2_0684_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2539_l2504_DUPLICATE_99f5_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2539_l2504_DUPLICATE_99f5_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
