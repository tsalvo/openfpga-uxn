-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity sub_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub_0CLK_bacf6a1d;
architecture arch of sub_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2336_c6_6b5a]
signal BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2336_c1_bff8]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2336_c2_8a05]
signal t8_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2336_c2_8a05]
signal n8_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2336_c2_8a05]
signal result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2336_c2_8a05]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2336_c2_8a05]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2336_c2_8a05]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2336_c2_8a05]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2336_c2_8a05]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l2337_c3_b04a[uxn_opcodes_h_l2337_c3_b04a]
signal printf_uxn_opcodes_h_l2337_c3_b04a_uxn_opcodes_h_l2337_c3_b04a_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2341_c11_2109]
signal BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2341_c7_84b6]
signal t8_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2341_c7_84b6]
signal n8_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2341_c7_84b6]
signal result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2341_c7_84b6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2341_c7_84b6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2341_c7_84b6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2341_c7_84b6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2341_c7_84b6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2344_c11_b204]
signal BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2344_c7_69e6]
signal t8_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2344_c7_69e6]
signal n8_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2344_c7_69e6]
signal result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2344_c7_69e6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2344_c7_69e6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2344_c7_69e6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2344_c7_69e6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2344_c7_69e6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2347_c11_d39a]
signal BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2347_c7_9f2c]
signal n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2347_c7_9f2c]
signal result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2347_c7_9f2c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2347_c7_9f2c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2347_c7_9f2c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2347_c7_9f2c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2347_c7_9f2c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2350_c30_a0ab]
signal sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_return_output : signed(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2353_c21_91a6]
signal BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2355_c11_43e0]
signal BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2355_c7_6260]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2355_c7_6260]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2355_c7_6260]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a
BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_left,
BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_right,
BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_return_output);

-- t8_MUX_uxn_opcodes_h_l2336_c2_8a05
t8_MUX_uxn_opcodes_h_l2336_c2_8a05 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2336_c2_8a05_cond,
t8_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue,
t8_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse,
t8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output);

-- n8_MUX_uxn_opcodes_h_l2336_c2_8a05
n8_MUX_uxn_opcodes_h_l2336_c2_8a05 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2336_c2_8a05_cond,
n8_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue,
n8_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse,
n8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05
result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_cond,
result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05
result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05
result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output);

-- printf_uxn_opcodes_h_l2337_c3_b04a_uxn_opcodes_h_l2337_c3_b04a
printf_uxn_opcodes_h_l2337_c3_b04a_uxn_opcodes_h_l2337_c3_b04a : entity work.printf_uxn_opcodes_h_l2337_c3_b04a_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2337_c3_b04a_uxn_opcodes_h_l2337_c3_b04a_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109
BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_left,
BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_right,
BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output);

-- t8_MUX_uxn_opcodes_h_l2341_c7_84b6
t8_MUX_uxn_opcodes_h_l2341_c7_84b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2341_c7_84b6_cond,
t8_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue,
t8_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse,
t8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output);

-- n8_MUX_uxn_opcodes_h_l2341_c7_84b6
n8_MUX_uxn_opcodes_h_l2341_c7_84b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2341_c7_84b6_cond,
n8_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue,
n8_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse,
n8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6
result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204
BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_left,
BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_right,
BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output);

-- t8_MUX_uxn_opcodes_h_l2344_c7_69e6
t8_MUX_uxn_opcodes_h_l2344_c7_69e6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2344_c7_69e6_cond,
t8_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue,
t8_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse,
t8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output);

-- n8_MUX_uxn_opcodes_h_l2344_c7_69e6
n8_MUX_uxn_opcodes_h_l2344_c7_69e6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2344_c7_69e6_cond,
n8_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue,
n8_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse,
n8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6
result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6
result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6
result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6
result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a
BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_left,
BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_right,
BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_return_output);

-- n8_MUX_uxn_opcodes_h_l2347_c7_9f2c
n8_MUX_uxn_opcodes_h_l2347_c7_9f2c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond,
n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue,
n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse,
n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c
result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c
result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c
result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c
result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab
sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_ins,
sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_x,
sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_y,
sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6
BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_left,
BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_right,
BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0
BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_left,
BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_right,
BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260
result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260
result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_return_output,
 t8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output,
 n8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output,
 t8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output,
 n8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output,
 t8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output,
 n8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_return_output,
 n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output,
 sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2338_c3_1aab : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2337_c3_b04a_uxn_opcodes_h_l2337_c3_b04a_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2342_c3_b1db : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2352_c3_7876 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_7eb8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_cfa3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_43b3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_0f74_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2344_l2347_l2341_l2355_DUPLICATE_240d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2344_l2347_DUPLICATE_0fc0_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2361_l2332_DUPLICATE_cfe4_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2352_c3_7876 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2352_c3_7876;
     VAR_sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2342_c3_b1db := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2342_c3_b1db;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_right := to_unsigned(3, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2338_c3_1aab := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2338_c3_1aab;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2336_c6_6b5a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2341_c11_2109] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_left;
     BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output := BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2355_c11_43e0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2350_c30_a0ab] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_ins;
     sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_x;
     sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_return_output := sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_cfa3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_cfa3_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2347_c11_d39a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2344_l2347_DUPLICATE_0fc0 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2344_l2347_DUPLICATE_0fc0_return_output := result.stack_address_sp_offset;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2353_c21_91a6] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_43b3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_43b3_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_0f74 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_0f74_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2344_l2347_l2341_l2355_DUPLICATE_240d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2344_l2347_l2341_l2355_DUPLICATE_240d_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_7eb8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_7eb8_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2344_c11_b204] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_left;
     BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output := BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2336_c2_8a05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2336_c2_8a05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c6_6b5a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2341_c7_84b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2341_c7_84b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_2109_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2344_c7_69e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2344_c7_69e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2344_c11_b204_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_d39a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_43e0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2353_c21_91a6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_0f74_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_0f74_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_0f74_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_0f74_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2344_l2347_l2341_l2355_DUPLICATE_240d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2344_l2347_l2341_l2355_DUPLICATE_240d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2344_l2347_l2341_l2355_DUPLICATE_240d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2344_l2347_l2341_l2355_DUPLICATE_240d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_cfa3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_cfa3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_cfa3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_cfa3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_43b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_43b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_43b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2344_l2336_l2341_l2355_DUPLICATE_43b3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2344_l2347_DUPLICATE_0fc0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2344_l2347_DUPLICATE_0fc0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_7eb8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_7eb8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_7eb8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2344_l2336_l2347_l2341_DUPLICATE_7eb8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2350_c30_a0ab_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2355_c7_6260] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_return_output;

     -- n8_MUX[uxn_opcodes_h_l2347_c7_9f2c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond;
     n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue;
     n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output := n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2336_c1_bff8] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2347_c7_9f2c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2347_c7_9f2c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;

     -- t8_MUX[uxn_opcodes_h_l2344_c7_69e6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2344_c7_69e6_cond <= VAR_t8_MUX_uxn_opcodes_h_l2344_c7_69e6_cond;
     t8_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue;
     t8_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output := t8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2355_c7_6260] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2347_c7_9f2c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2355_c7_6260] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2337_c3_b04a_uxn_opcodes_h_l2337_c3_b04a_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2336_c1_bff8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_6260_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2355_c7_6260_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_6260_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2347_c7_9f2c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;

     -- printf_uxn_opcodes_h_l2337_c3_b04a[uxn_opcodes_h_l2337_c3_b04a] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2337_c3_b04a_uxn_opcodes_h_l2337_c3_b04a_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2337_c3_b04a_uxn_opcodes_h_l2337_c3_b04a_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2344_c7_69e6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;

     -- n8_MUX[uxn_opcodes_h_l2344_c7_69e6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2344_c7_69e6_cond <= VAR_n8_MUX_uxn_opcodes_h_l2344_c7_69e6_cond;
     n8_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue;
     n8_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output := n8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;

     -- t8_MUX[uxn_opcodes_h_l2341_c7_84b6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2341_c7_84b6_cond <= VAR_t8_MUX_uxn_opcodes_h_l2341_c7_84b6_cond;
     t8_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue;
     t8_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output := t8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2344_c7_69e6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2347_c7_9f2c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2347_c7_9f2c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2344_c7_69e6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_9f2c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;
     -- t8_MUX[uxn_opcodes_h_l2336_c2_8a05] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2336_c2_8a05_cond <= VAR_t8_MUX_uxn_opcodes_h_l2336_c2_8a05_cond;
     t8_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue;
     t8_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output := t8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2344_c7_69e6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;

     -- n8_MUX[uxn_opcodes_h_l2341_c7_84b6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2341_c7_84b6_cond <= VAR_n8_MUX_uxn_opcodes_h_l2341_c7_84b6_cond;
     n8_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue;
     n8_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output := n8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2341_c7_84b6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2344_c7_69e6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2344_c7_69e6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2341_c7_84b6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2341_c7_84b6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2344_c7_69e6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2341_c7_84b6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2336_c2_8a05] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2341_c7_84b6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;

     -- n8_MUX[uxn_opcodes_h_l2336_c2_8a05] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2336_c2_8a05_cond <= VAR_n8_MUX_uxn_opcodes_h_l2336_c2_8a05_cond;
     n8_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue;
     n8_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output := n8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2336_c2_8a05] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output := result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2341_c7_84b6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2336_c2_8a05] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_84b6_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2336_c2_8a05] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2336_c2_8a05] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2336_c2_8a05] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2361_l2332_DUPLICATE_cfe4 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2361_l2332_DUPLICATE_cfe4_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c2_8a05_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2361_l2332_DUPLICATE_cfe4_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2361_l2332_DUPLICATE_cfe4_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
