-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity equ2_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end equ2_0CLK_85d5529e;
architecture arch of equ2_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1093_c6_799e]
signal BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1093_c2_3a62]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1093_c2_3a62]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1093_c2_3a62]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1093_c2_3a62]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1093_c2_3a62]
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1093_c2_3a62]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1093_c2_3a62]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1093_c2_3a62]
signal n16_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1093_c2_3a62]
signal t16_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1101_c11_d9e1]
signal BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1101_c7_f2fa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1101_c7_f2fa]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1101_c7_f2fa]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1101_c7_f2fa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1101_c7_f2fa]
signal result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1101_c7_f2fa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1101_c7_f2fa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1101_c7_f2fa]
signal n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1101_c7_f2fa]
signal t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1104_c11_07dd]
signal BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1104_c7_62c6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1104_c7_62c6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1104_c7_62c6]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1104_c7_62c6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1104_c7_62c6]
signal result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1104_c7_62c6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1104_c7_62c6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1104_c7_62c6]
signal n16_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1104_c7_62c6]
signal t16_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1108_c30_f2a1]
signal sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1110_c11_7531]
signal BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1110_c7_fa9b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1110_c7_fa9b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1110_c7_fa9b]
signal result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1110_c7_fa9b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1110_c7_fa9b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l1110_c7_fa9b]
signal n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1115_c21_6048]
signal BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_left : unsigned(15 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_right : unsigned(15 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1115_c21_afc7]
signal MUX_uxn_opcodes_h_l1115_c21_afc7_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1115_c21_afc7_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1115_c21_afc7_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1115_c21_afc7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1117_c11_f86a]
signal BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1117_c7_57f6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1117_c7_57f6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_stack_operation_16bit := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e
BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_left,
BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_right,
BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62
result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62
result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_cond,
result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output);

-- n16_MUX_uxn_opcodes_h_l1093_c2_3a62
n16_MUX_uxn_opcodes_h_l1093_c2_3a62 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1093_c2_3a62_cond,
n16_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue,
n16_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse,
n16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output);

-- t16_MUX_uxn_opcodes_h_l1093_c2_3a62
t16_MUX_uxn_opcodes_h_l1093_c2_3a62 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1093_c2_3a62_cond,
t16_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue,
t16_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse,
t16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1
BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_left,
BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_right,
BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa
result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa
result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa
result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond,
result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa
result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa
result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output);

-- n16_MUX_uxn_opcodes_h_l1101_c7_f2fa
n16_MUX_uxn_opcodes_h_l1101_c7_f2fa : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond,
n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue,
n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse,
n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output);

-- t16_MUX_uxn_opcodes_h_l1101_c7_f2fa
t16_MUX_uxn_opcodes_h_l1101_c7_f2fa : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond,
t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue,
t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse,
t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd
BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_left,
BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_right,
BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6
result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6
result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6
result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_cond,
result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6
result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6
result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output);

-- n16_MUX_uxn_opcodes_h_l1104_c7_62c6
n16_MUX_uxn_opcodes_h_l1104_c7_62c6 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1104_c7_62c6_cond,
n16_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue,
n16_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse,
n16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output);

-- t16_MUX_uxn_opcodes_h_l1104_c7_62c6
t16_MUX_uxn_opcodes_h_l1104_c7_62c6 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1104_c7_62c6_cond,
t16_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue,
t16_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse,
t16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1
sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_ins,
sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_x,
sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_y,
sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531
BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_left,
BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_right,
BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b
result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b
result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b
result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b
result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output);

-- n16_MUX_uxn_opcodes_h_l1110_c7_fa9b
n16_MUX_uxn_opcodes_h_l1110_c7_fa9b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond,
n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue,
n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse,
n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048
BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048 : entity work.BIN_OP_EQ_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_left,
BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_right,
BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_return_output);

-- MUX_uxn_opcodes_h_l1115_c21_afc7
MUX_uxn_opcodes_h_l1115_c21_afc7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1115_c21_afc7_cond,
MUX_uxn_opcodes_h_l1115_c21_afc7_iftrue,
MUX_uxn_opcodes_h_l1115_c21_afc7_iffalse,
MUX_uxn_opcodes_h_l1115_c21_afc7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a
BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_left,
BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_right,
BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6
result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6
result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
 n16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
 t16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output,
 n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output,
 t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output,
 n16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output,
 t16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output,
 sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output,
 n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_return_output,
 MUX_uxn_opcodes_h_l1115_c21_afc7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1098_c3_2dc4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1093_c2_3a62_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1102_c3_855c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1104_c7_62c6_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1114_c3_8557 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1115_c21_afc7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1115_c21_afc7_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1115_c21_afc7_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1115_c21_afc7_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1101_l1110_l1093_DUPLICATE_afc9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1101_l1110_l1093_l1104_DUPLICATE_45d5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1101_l1093_l1104_DUPLICATE_8bca_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1117_l1101_l1093_l1104_DUPLICATE_717f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1101_l1104_DUPLICATE_5d95_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1117_l1101_l1110_l1104_DUPLICATE_bda7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1110_l1104_DUPLICATE_d189_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1122_l1089_DUPLICATE_dff6_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_y := resize(to_signed(-3, 3), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1102_c3_855c := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1102_c3_855c;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1114_c3_8557 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1114_c3_8557;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1098_c3_2dc4 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1098_c3_2dc4;
     VAR_MUX_uxn_opcodes_h_l1115_c21_afc7_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1115_c21_afc7_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_left := VAR_previous_stack_read;
     VAR_n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_right := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse := t16;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1101_l1093_l1104_DUPLICATE_8bca LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1101_l1093_l1104_DUPLICATE_8bca_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1104_c11_07dd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_left;
     BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output := BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1101_l1110_l1093_l1104_DUPLICATE_45d5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1101_l1110_l1093_l1104_DUPLICATE_45d5_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1093_c6_799e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1110_c11_7531] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_left;
     BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_return_output := BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1115_c21_6048] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_left;
     BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_return_output := BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1101_c11_d9e1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1117_c11_f86a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1101_l1104_DUPLICATE_5d95 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1101_l1104_DUPLICATE_5d95_return_output := result.is_stack_operation_16bit;

     -- sp_relative_shift[uxn_opcodes_h_l1108_c30_f2a1] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_ins;
     sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_x;
     sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_return_output := sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1101_l1110_l1093_DUPLICATE_afc9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1101_l1110_l1093_DUPLICATE_afc9_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1110_l1104_DUPLICATE_d189 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1110_l1104_DUPLICATE_d189_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1117_l1101_l1110_l1104_DUPLICATE_bda7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1117_l1101_l1110_l1104_DUPLICATE_bda7_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1117_l1101_l1093_l1104_DUPLICATE_717f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1117_l1101_l1093_l1104_DUPLICATE_717f_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_n16_MUX_uxn_opcodes_h_l1093_c2_3a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1093_c2_3a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c6_799e_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1101_c11_d9e1_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1104_c7_62c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1104_c7_62c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1104_c11_07dd_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1110_c11_7531_return_output;
     VAR_MUX_uxn_opcodes_h_l1115_c21_afc7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c21_6048_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1117_c11_f86a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1101_l1093_l1104_DUPLICATE_8bca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1101_l1093_l1104_DUPLICATE_8bca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1101_l1093_l1104_DUPLICATE_8bca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1117_l1101_l1110_l1104_DUPLICATE_bda7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1117_l1101_l1110_l1104_DUPLICATE_bda7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1117_l1101_l1110_l1104_DUPLICATE_bda7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1117_l1101_l1110_l1104_DUPLICATE_bda7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1101_l1110_l1093_DUPLICATE_afc9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1101_l1110_l1093_DUPLICATE_afc9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1101_l1110_l1093_DUPLICATE_afc9_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1101_l1104_DUPLICATE_5d95_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1101_l1104_DUPLICATE_5d95_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1117_l1101_l1093_l1104_DUPLICATE_717f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1117_l1101_l1093_l1104_DUPLICATE_717f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1117_l1101_l1093_l1104_DUPLICATE_717f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1117_l1101_l1093_l1104_DUPLICATE_717f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1110_l1104_DUPLICATE_d189_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1110_l1104_DUPLICATE_d189_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1101_l1110_l1093_l1104_DUPLICATE_45d5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1101_l1110_l1093_l1104_DUPLICATE_45d5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1101_l1110_l1093_l1104_DUPLICATE_45d5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1101_l1110_l1093_l1104_DUPLICATE_45d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1108_c30_f2a1_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1104_c7_62c6] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;

     -- MUX[uxn_opcodes_h_l1115_c21_afc7] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1115_c21_afc7_cond <= VAR_MUX_uxn_opcodes_h_l1115_c21_afc7_cond;
     MUX_uxn_opcodes_h_l1115_c21_afc7_iftrue <= VAR_MUX_uxn_opcodes_h_l1115_c21_afc7_iftrue;
     MUX_uxn_opcodes_h_l1115_c21_afc7_iffalse <= VAR_MUX_uxn_opcodes_h_l1115_c21_afc7_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1115_c21_afc7_return_output := MUX_uxn_opcodes_h_l1115_c21_afc7_return_output;

     -- t16_MUX[uxn_opcodes_h_l1104_c7_62c6] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1104_c7_62c6_cond <= VAR_t16_MUX_uxn_opcodes_h_l1104_c7_62c6_cond;
     t16_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue;
     t16_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output := t16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1117_c7_57f6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1117_c7_57f6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1104_c7_62c6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1110_c7_fa9b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1110_c7_fa9b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output;

     -- n16_MUX[uxn_opcodes_h_l1110_c7_fa9b] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond <= VAR_n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond;
     n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue;
     n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output := n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue := VAR_MUX_uxn_opcodes_h_l1115_c21_afc7_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1117_c7_57f6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;
     -- n16_MUX[uxn_opcodes_h_l1104_c7_62c6] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1104_c7_62c6_cond <= VAR_n16_MUX_uxn_opcodes_h_l1104_c7_62c6_cond;
     n16_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue;
     n16_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output := n16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1101_c7_f2fa] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1110_c7_fa9b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output;

     -- t16_MUX[uxn_opcodes_h_l1101_c7_f2fa] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond <= VAR_t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond;
     t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue;
     t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output := t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1104_c7_62c6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1104_c7_62c6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1110_c7_fa9b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1110_c7_fa9b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1101_c7_f2fa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1110_c7_fa9b_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1093_c2_3a62] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1104_c7_62c6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1104_c7_62c6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output := result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1101_c7_f2fa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;

     -- t16_MUX[uxn_opcodes_h_l1093_c2_3a62] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1093_c2_3a62_cond <= VAR_t16_MUX_uxn_opcodes_h_l1093_c2_3a62_cond;
     t16_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue;
     t16_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output := t16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1101_c7_f2fa] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;

     -- n16_MUX[uxn_opcodes_h_l1101_c7_f2fa] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond <= VAR_n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond;
     n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue;
     n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output := n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1093_c2_3a62] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1104_c7_62c6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1104_c7_62c6_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1101_c7_f2fa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;

     -- n16_MUX[uxn_opcodes_h_l1093_c2_3a62] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1093_c2_3a62_cond <= VAR_n16_MUX_uxn_opcodes_h_l1093_c2_3a62_cond;
     n16_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue;
     n16_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output := n16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1093_c2_3a62] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1101_c7_f2fa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1101_c7_f2fa] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output := result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1093_c2_3a62] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1101_c7_f2fa_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1093_c2_3a62] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1093_c2_3a62] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output := result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1093_c2_3a62] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1122_l1089_DUPLICATE_dff6 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1122_l1089_DUPLICATE_dff6_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c2_3a62_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1122_l1089_DUPLICATE_dff6_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1122_l1089_DUPLICATE_dff6_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
