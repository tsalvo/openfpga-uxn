-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity neq_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_226c8821;
architecture arch of neq_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1242_c6_1d50]
signal BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1242_c2_62e5]
signal n8_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1242_c2_62e5]
signal t8_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1242_c2_62e5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1242_c2_62e5]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1242_c2_62e5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1242_c2_62e5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1242_c2_62e5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1242_c2_62e5]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1242_c2_62e5]
signal result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1242_c2_62e5]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1242_c2_62e5]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1255_c11_6c8a]
signal BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1255_c7_8528]
signal n8_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1255_c7_8528]
signal t8_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1255_c7_8528]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1255_c7_8528]
signal result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1255_c7_8528]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1255_c7_8528]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1255_c7_8528]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1258_c11_f858]
signal BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1258_c7_62a4]
signal n8_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1258_c7_62a4]
signal t8_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1258_c7_62a4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1258_c7_62a4]
signal result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1258_c7_62a4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1258_c7_62a4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1258_c7_62a4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1261_c11_dab1]
signal BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1261_c7_43b3]
signal n8_MUX_uxn_opcodes_h_l1261_c7_43b3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1261_c7_43b3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1261_c7_43b3]
signal result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1261_c7_43b3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1261_c7_43b3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1261_c7_43b3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1263_c30_2901]
signal sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1266_c21_2aa0]
signal BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1266_c21_abdc]
signal MUX_uxn_opcodes_h_l1266_c21_abdc_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1266_c21_abdc_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1266_c21_abdc_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1266_c21_abdc_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_ee25( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_vram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50
BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_left,
BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_right,
BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output);

-- n8_MUX_uxn_opcodes_h_l1242_c2_62e5
n8_MUX_uxn_opcodes_h_l1242_c2_62e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1242_c2_62e5_cond,
n8_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue,
n8_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse,
n8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output);

-- t8_MUX_uxn_opcodes_h_l1242_c2_62e5
t8_MUX_uxn_opcodes_h_l1242_c2_62e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1242_c2_62e5_cond,
t8_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue,
t8_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse,
t8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a
BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_left,
BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_right,
BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_return_output);

-- n8_MUX_uxn_opcodes_h_l1255_c7_8528
n8_MUX_uxn_opcodes_h_l1255_c7_8528 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1255_c7_8528_cond,
n8_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue,
n8_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse,
n8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output);

-- t8_MUX_uxn_opcodes_h_l1255_c7_8528
t8_MUX_uxn_opcodes_h_l1255_c7_8528 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1255_c7_8528_cond,
t8_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue,
t8_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse,
t8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_cond,
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858
BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_left,
BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_right,
BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_return_output);

-- n8_MUX_uxn_opcodes_h_l1258_c7_62a4
n8_MUX_uxn_opcodes_h_l1258_c7_62a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1258_c7_62a4_cond,
n8_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue,
n8_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse,
n8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output);

-- t8_MUX_uxn_opcodes_h_l1258_c7_62a4
t8_MUX_uxn_opcodes_h_l1258_c7_62a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1258_c7_62a4_cond,
t8_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue,
t8_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse,
t8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1
BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_left,
BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_right,
BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_return_output);

-- n8_MUX_uxn_opcodes_h_l1261_c7_43b3
n8_MUX_uxn_opcodes_h_l1261_c7_43b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1261_c7_43b3_cond,
n8_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue,
n8_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse,
n8_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_cond,
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1263_c30_2901
sp_relative_shift_uxn_opcodes_h_l1263_c30_2901 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_ins,
sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_x,
sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_y,
sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0
BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_left,
BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_right,
BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_return_output);

-- MUX_uxn_opcodes_h_l1266_c21_abdc
MUX_uxn_opcodes_h_l1266_c21_abdc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1266_c21_abdc_cond,
MUX_uxn_opcodes_h_l1266_c21_abdc_iftrue,
MUX_uxn_opcodes_h_l1266_c21_abdc_iffalse,
MUX_uxn_opcodes_h_l1266_c21_abdc_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output,
 n8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
 t8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_return_output,
 n8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output,
 t8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_return_output,
 n8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output,
 t8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_return_output,
 n8_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output,
 sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_return_output,
 MUX_uxn_opcodes_h_l1266_c21_abdc_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1247_c3_5482 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1252_c3_5be4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1256_c3_8db0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1261_c7_43b3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1265_c3_f034 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1266_c21_abdc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1266_c21_abdc_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1266_c21_abdc_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1266_c21_abdc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1258_l1242_l1261_l1255_DUPLICATE_f6e7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_2ef9_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_a81e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_d174_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_a315_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l1270_l1238_DUPLICATE_5654_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1247_c3_5482 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1247_c3_5482;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1265_c3_f034 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1265_c3_f034;
     VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_right := to_unsigned(3, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1256_c3_8db0 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1256_c3_8db0;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_right := to_unsigned(2, 2);
     VAR_MUX_uxn_opcodes_h_l1266_c21_abdc_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1252_c3_5be4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1252_c3_5be4;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1266_c21_abdc_iffalse := resize(to_unsigned(1, 1), 8);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_2ef9 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_2ef9_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1266_c21_2aa0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_a315 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_a315_return_output := result.stack_address_sp_offset;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1242_c2_62e5_return_output := result.is_ram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1242_c2_62e5_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l1263_c30_2901] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_ins;
     sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_x;
     sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_return_output := sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1255_c11_6c8a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_d174 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_d174_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1258_c11_f858] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_left;
     BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_return_output := BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1242_c2_62e5_return_output := result.is_vram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1242_c2_62e5_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1258_l1242_l1261_l1255_DUPLICATE_f6e7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1258_l1242_l1261_l1255_DUPLICATE_f6e7_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_a81e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_a81e_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1242_c6_1d50] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_left;
     BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output := BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1261_c11_dab1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1242_c2_62e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1242_c2_62e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_1d50_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1255_c7_8528_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1255_c7_8528_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_6c8a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1258_c7_62a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1258_c7_62a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_f858_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1261_c7_43b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_dab1_return_output;
     VAR_MUX_uxn_opcodes_h_l1266_c21_abdc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_2aa0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_2ef9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_2ef9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_2ef9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_d174_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_d174_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_d174_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_a81e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_a81e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1258_l1261_l1255_DUPLICATE_a81e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_a315_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_a315_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1258_l1242_l1261_l1255_DUPLICATE_f6e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1258_l1242_l1261_l1255_DUPLICATE_f6e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1258_l1242_l1261_l1255_DUPLICATE_f6e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1258_l1242_l1261_l1255_DUPLICATE_f6e7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1242_c2_62e5_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1242_c2_62e5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1242_c2_62e5_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1242_c2_62e5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_2901_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1261_c7_43b3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1261_c7_43b3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1261_c7_43b3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1261_c7_43b3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output;

     -- MUX[uxn_opcodes_h_l1266_c21_abdc] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1266_c21_abdc_cond <= VAR_MUX_uxn_opcodes_h_l1266_c21_abdc_cond;
     MUX_uxn_opcodes_h_l1266_c21_abdc_iftrue <= VAR_MUX_uxn_opcodes_h_l1266_c21_abdc_iftrue;
     MUX_uxn_opcodes_h_l1266_c21_abdc_iffalse <= VAR_MUX_uxn_opcodes_h_l1266_c21_abdc_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1266_c21_abdc_return_output := MUX_uxn_opcodes_h_l1266_c21_abdc_return_output;

     -- t8_MUX[uxn_opcodes_h_l1258_c7_62a4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1258_c7_62a4_cond <= VAR_t8_MUX_uxn_opcodes_h_l1258_c7_62a4_cond;
     t8_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue;
     t8_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output := t8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1261_c7_43b3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1261_c7_43b3_cond <= VAR_n8_MUX_uxn_opcodes_h_l1261_c7_43b3_cond;
     n8_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue;
     n8_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output := n8_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue := VAR_MUX_uxn_opcodes_h_l1266_c21_abdc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;
     -- t8_MUX[uxn_opcodes_h_l1255_c7_8528] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1255_c7_8528_cond <= VAR_t8_MUX_uxn_opcodes_h_l1255_c7_8528_cond;
     t8_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue;
     t8_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output := t8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1258_c7_62a4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1258_c7_62a4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1258_c7_62a4_cond <= VAR_n8_MUX_uxn_opcodes_h_l1258_c7_62a4_cond;
     n8_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue;
     n8_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output := n8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1258_c7_62a4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1261_c7_43b3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output := result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1258_c7_62a4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1258_c7_62a4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_43b3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;
     -- t8_MUX[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1242_c2_62e5_cond <= VAR_t8_MUX_uxn_opcodes_h_l1242_c2_62e5_cond;
     t8_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue;
     t8_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output := t8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output;

     -- n8_MUX[uxn_opcodes_h_l1255_c7_8528] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1255_c7_8528_cond <= VAR_n8_MUX_uxn_opcodes_h_l1255_c7_8528_cond;
     n8_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue;
     n8_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output := n8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1255_c7_8528] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1255_c7_8528] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1255_c7_8528] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1255_c7_8528] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1258_c7_62a4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_62a4_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output;
     -- n8_MUX[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1242_c2_62e5_cond <= VAR_n8_MUX_uxn_opcodes_h_l1242_c2_62e5_cond;
     n8_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue;
     n8_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output := n8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1255_c7_8528] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_return_output := result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_8528_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1242_c2_62e5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l1270_l1238_DUPLICATE_5654 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l1270_l1238_DUPLICATE_5654_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_ee25(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_62e5_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l1270_l1238_DUPLICATE_5654_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l1270_l1238_DUPLICATE_5654_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
