-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity lth_0CLK_441a128d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lth_0CLK_441a128d;
architecture arch of lth_0CLK_441a128d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1890_c6_e427]
signal BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1890_c2_3eda]
signal n8_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1890_c2_3eda]
signal t8_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1890_c2_3eda]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1890_c2_3eda]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1890_c2_3eda]
signal result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1890_c2_3eda]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1890_c2_3eda]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1890_c2_3eda]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1890_c2_3eda]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1890_c2_3eda]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1890_c2_3eda]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1903_c11_c4c5]
signal BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1903_c7_738d]
signal n8_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1903_c7_738d]
signal t8_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1903_c7_738d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1903_c7_738d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1903_c7_738d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1903_c7_738d]
signal result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1903_c7_738d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1906_c11_11e1]
signal BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1906_c7_987f]
signal n8_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1906_c7_987f]
signal t8_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1906_c7_987f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1906_c7_987f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1906_c7_987f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1906_c7_987f]
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1906_c7_987f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1909_c11_7b61]
signal BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1909_c7_1f6b]
signal n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1909_c7_1f6b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1909_c7_1f6b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1909_c7_1f6b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1909_c7_1f6b]
signal result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1909_c7_1f6b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1911_c30_8cdf]
signal sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_return_output : signed(3 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l1914_c21_9ab1]
signal BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1914_c21_8819]
signal MUX_uxn_opcodes_h_l1914_c21_8819_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1914_c21_8819_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1914_c21_8819_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1914_c21_8819_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a6df( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_vram_write := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427
BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_left,
BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_right,
BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output);

-- n8_MUX_uxn_opcodes_h_l1890_c2_3eda
n8_MUX_uxn_opcodes_h_l1890_c2_3eda : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1890_c2_3eda_cond,
n8_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue,
n8_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse,
n8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output);

-- t8_MUX_uxn_opcodes_h_l1890_c2_3eda
t8_MUX_uxn_opcodes_h_l1890_c2_3eda : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1890_c2_3eda_cond,
t8_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue,
t8_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse,
t8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda
result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda
result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_cond,
result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda
result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda
result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda
result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda
result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda
result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5
BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_left,
BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_right,
BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_return_output);

-- n8_MUX_uxn_opcodes_h_l1903_c7_738d
n8_MUX_uxn_opcodes_h_l1903_c7_738d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1903_c7_738d_cond,
n8_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue,
n8_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse,
n8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output);

-- t8_MUX_uxn_opcodes_h_l1903_c7_738d
t8_MUX_uxn_opcodes_h_l1903_c7_738d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1903_c7_738d_cond,
t8_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue,
t8_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse,
t8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d
result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d
result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d
result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1
BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_left,
BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_right,
BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_return_output);

-- n8_MUX_uxn_opcodes_h_l1906_c7_987f
n8_MUX_uxn_opcodes_h_l1906_c7_987f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1906_c7_987f_cond,
n8_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue,
n8_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse,
n8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output);

-- t8_MUX_uxn_opcodes_h_l1906_c7_987f
t8_MUX_uxn_opcodes_h_l1906_c7_987f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1906_c7_987f_cond,
t8_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue,
t8_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse,
t8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f
result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61
BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_left,
BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_right,
BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_return_output);

-- n8_MUX_uxn_opcodes_h_l1909_c7_1f6b
n8_MUX_uxn_opcodes_h_l1909_c7_1f6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond,
n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue,
n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse,
n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b
result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b
result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b
result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf
sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_ins,
sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_x,
sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_y,
sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1
BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1 : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_380ecc95 port map (
BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_left,
BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_right,
BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_return_output);

-- MUX_uxn_opcodes_h_l1914_c21_8819
MUX_uxn_opcodes_h_l1914_c21_8819 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1914_c21_8819_cond,
MUX_uxn_opcodes_h_l1914_c21_8819_iftrue,
MUX_uxn_opcodes_h_l1914_c21_8819_iffalse,
MUX_uxn_opcodes_h_l1914_c21_8819_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output,
 n8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
 t8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_return_output,
 n8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output,
 t8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_return_output,
 n8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output,
 t8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_return_output,
 n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output,
 sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_return_output,
 BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_return_output,
 MUX_uxn_opcodes_h_l1914_c21_8819_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1895_c3_d46d : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1900_c3_cee1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1904_c3_aabb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1913_c3_1c5f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1914_c21_8819_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1914_c21_8819_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1914_c21_8819_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1914_c21_8819_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1890_l1909_l1903_l1906_DUPLICATE_84b0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_c0fb_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_b33c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_6ab5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1909_l1906_DUPLICATE_4aac_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1918_l1886_DUPLICATE_346b_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1914_c21_8819_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_right := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1904_c3_aabb := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1904_c3_aabb;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1913_c3_1c5f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1913_c3_1c5f;
     VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1900_c3_cee1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1900_c3_cee1;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_y := resize(to_signed(-1, 2), 4);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1895_c3_d46d := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1895_c3_d46d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1914_c21_8819_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse := t8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1909_l1906_DUPLICATE_4aac LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1909_l1906_DUPLICATE_4aac_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_c0fb LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_c0fb_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l1911_c30_8cdf] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_ins;
     sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_x;
     sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_return_output := sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_return_output;

     -- BIN_OP_LT[uxn_opcodes_h_l1914_c21_9ab1] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_left;
     BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_return_output := BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1890_c2_3eda_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_b33c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_b33c_return_output := result.is_opc_done;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1890_c2_3eda_return_output := result.is_ram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1890_c2_3eda_return_output := result.is_pc_updated;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1890_c2_3eda_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_6ab5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_6ab5_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1903_c11_c4c5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1890_l1909_l1903_l1906_DUPLICATE_84b0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1890_l1909_l1903_l1906_DUPLICATE_84b0_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1906_c11_11e1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1909_c11_7b61] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_left;
     BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_return_output := BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1890_c6_e427] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_left;
     BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output := BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1890_c2_3eda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1890_c2_3eda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_e427_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1903_c7_738d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1903_c7_738d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_c4c5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1906_c7_987f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1906_c7_987f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_11e1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_7b61_return_output;
     VAR_MUX_uxn_opcodes_h_l1914_c21_8819_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_9ab1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_c0fb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_c0fb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_c0fb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_b33c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_b33c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_b33c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_6ab5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_6ab5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1909_l1903_l1906_DUPLICATE_6ab5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1909_l1906_DUPLICATE_4aac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1909_l1906_DUPLICATE_4aac_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1890_l1909_l1903_l1906_DUPLICATE_84b0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1890_l1909_l1903_l1906_DUPLICATE_84b0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1890_l1909_l1903_l1906_DUPLICATE_84b0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1890_l1909_l1903_l1906_DUPLICATE_84b0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1890_c2_3eda_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1890_c2_3eda_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1890_c2_3eda_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1890_c2_3eda_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_8cdf_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1909_c7_1f6b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1906_c7_987f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1906_c7_987f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1906_c7_987f_cond;
     t8_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue;
     t8_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output := t8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1909_c7_1f6b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output;

     -- MUX[uxn_opcodes_h_l1914_c21_8819] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1914_c21_8819_cond <= VAR_MUX_uxn_opcodes_h_l1914_c21_8819_cond;
     MUX_uxn_opcodes_h_l1914_c21_8819_iftrue <= VAR_MUX_uxn_opcodes_h_l1914_c21_8819_iftrue;
     MUX_uxn_opcodes_h_l1914_c21_8819_iffalse <= VAR_MUX_uxn_opcodes_h_l1914_c21_8819_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1914_c21_8819_return_output := MUX_uxn_opcodes_h_l1914_c21_8819_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output;

     -- n8_MUX[uxn_opcodes_h_l1909_c7_1f6b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond;
     n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue;
     n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output := n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1909_c7_1f6b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1909_c7_1f6b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue := VAR_MUX_uxn_opcodes_h_l1914_c21_8819_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1906_c7_987f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1906_c7_987f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1909_c7_1f6b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output;

     -- n8_MUX[uxn_opcodes_h_l1906_c7_987f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1906_c7_987f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1906_c7_987f_cond;
     n8_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue;
     n8_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output := n8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1903_c7_738d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1903_c7_738d_cond <= VAR_t8_MUX_uxn_opcodes_h_l1903_c7_738d_cond;
     t8_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue;
     t8_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output := t8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1906_c7_987f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1906_c7_987f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_1f6b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;
     -- n8_MUX[uxn_opcodes_h_l1903_c7_738d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1903_c7_738d_cond <= VAR_n8_MUX_uxn_opcodes_h_l1903_c7_738d_cond;
     n8_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue;
     n8_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output := n8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1903_c7_738d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1903_c7_738d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1906_c7_987f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1890_c2_3eda_cond <= VAR_t8_MUX_uxn_opcodes_h_l1890_c2_3eda_cond;
     t8_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue;
     t8_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output := t8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1903_c7_738d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1903_c7_738d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_987f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output;

     -- n8_MUX[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1890_c2_3eda_cond <= VAR_n8_MUX_uxn_opcodes_h_l1890_c2_3eda_cond;
     n8_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue;
     n8_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output := n8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1903_c7_738d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_738d_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1890_c2_3eda] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output := result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1918_l1886_DUPLICATE_346b LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1918_l1886_DUPLICATE_346b_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a6df(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_3eda_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1918_l1886_DUPLICATE_346b_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1918_l1886_DUPLICATE_346b_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
