-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity ora_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ora_0CLK_bacf6a1d;
architecture arch of ora_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l956_c6_d13e]
signal BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l956_c1_02c9]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l956_c2_cbea]
signal n8_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l956_c2_cbea]
signal t8_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l956_c2_cbea]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l956_c2_cbea]
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l956_c2_cbea]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l956_c2_cbea]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l956_c2_cbea]
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l956_c2_cbea]
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l957_c3_0a25[uxn_opcodes_h_l957_c3_0a25]
signal printf_uxn_opcodes_h_l957_c3_0a25_uxn_opcodes_h_l957_c3_0a25_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l961_c11_353a]
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l961_c7_fc74]
signal n8_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l961_c7_fc74]
signal t8_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l961_c7_fc74]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l961_c7_fc74]
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l961_c7_fc74]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l961_c7_fc74]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l961_c7_fc74]
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l961_c7_fc74]
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l964_c11_9b1e]
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l964_c7_5cff]
signal n8_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l964_c7_5cff]
signal t8_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l964_c7_5cff]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l964_c7_5cff]
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l964_c7_5cff]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l964_c7_5cff]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l964_c7_5cff]
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l964_c7_5cff]
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l967_c11_eb1a]
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l967_c7_805f]
signal n8_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l967_c7_805f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l967_c7_805f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l967_c7_805f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l967_c7_805f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l967_c7_805f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l967_c7_805f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l967_c7_805f]
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l970_c30_f07a]
signal sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l973_c21_010e]
signal BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_left : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_right : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l975_c11_661d]
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l975_c7_df82]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l975_c7_df82]
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l975_c7_df82]
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_4e73( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e
BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_left,
BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_right,
BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_return_output);

-- n8_MUX_uxn_opcodes_h_l956_c2_cbea
n8_MUX_uxn_opcodes_h_l956_c2_cbea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l956_c2_cbea_cond,
n8_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue,
n8_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse,
n8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output);

-- t8_MUX_uxn_opcodes_h_l956_c2_cbea
t8_MUX_uxn_opcodes_h_l956_c2_cbea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l956_c2_cbea_cond,
t8_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue,
t8_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse,
t8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea
result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_cond,
result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_return_output);

-- printf_uxn_opcodes_h_l957_c3_0a25_uxn_opcodes_h_l957_c3_0a25
printf_uxn_opcodes_h_l957_c3_0a25_uxn_opcodes_h_l957_c3_0a25 : entity work.printf_uxn_opcodes_h_l957_c3_0a25_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l957_c3_0a25_uxn_opcodes_h_l957_c3_0a25_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a
BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_left,
BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_right,
BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output);

-- n8_MUX_uxn_opcodes_h_l961_c7_fc74
n8_MUX_uxn_opcodes_h_l961_c7_fc74 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l961_c7_fc74_cond,
n8_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue,
n8_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse,
n8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output);

-- t8_MUX_uxn_opcodes_h_l961_c7_fc74
t8_MUX_uxn_opcodes_h_l961_c7_fc74 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l961_c7_fc74_cond,
t8_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue,
t8_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse,
t8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74
result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_cond,
result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e
BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_left,
BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_right,
BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output);

-- n8_MUX_uxn_opcodes_h_l964_c7_5cff
n8_MUX_uxn_opcodes_h_l964_c7_5cff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l964_c7_5cff_cond,
n8_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue,
n8_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse,
n8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output);

-- t8_MUX_uxn_opcodes_h_l964_c7_5cff
t8_MUX_uxn_opcodes_h_l964_c7_5cff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l964_c7_5cff_cond,
t8_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue,
t8_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse,
t8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff
result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_cond,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a
BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_left,
BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_right,
BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_return_output);

-- n8_MUX_uxn_opcodes_h_l967_c7_805f
n8_MUX_uxn_opcodes_h_l967_c7_805f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l967_c7_805f_cond,
n8_MUX_uxn_opcodes_h_l967_c7_805f_iftrue,
n8_MUX_uxn_opcodes_h_l967_c7_805f_iffalse,
n8_MUX_uxn_opcodes_h_l967_c7_805f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f
result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_cond,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_return_output);

-- sp_relative_shift_uxn_opcodes_h_l970_c30_f07a
sp_relative_shift_uxn_opcodes_h_l970_c30_f07a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_ins,
sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_x,
sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_y,
sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l973_c21_010e
BIN_OP_OR_uxn_opcodes_h_l973_c21_010e : entity work.BIN_OP_OR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_left,
BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_right,
BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d
BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_left,
BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_right,
BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_return_output,
 n8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output,
 t8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output,
 n8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output,
 t8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output,
 n8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output,
 t8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_return_output,
 n8_MUX_uxn_opcodes_h_l967_c7_805f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_return_output,
 sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_return_output,
 BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_c1ba : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l957_c3_0a25_uxn_opcodes_h_l957_c3_0a25_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_18e8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_805f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_8d5b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_bd47_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_2a6c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_75f2_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_6a03_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l967_l961_l975_l964_DUPLICATE_c598_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l967_l964_DUPLICATE_60df_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l952_l981_DUPLICATE_8b0f_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_8d5b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l972_c3_8d5b;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_18e8 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l962_c3_18e8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_c1ba := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l958_c3_c1ba;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_805f_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_805f_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l970_c30_f07a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_ins;
     sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_x;
     sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_return_output := sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_bd47 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_bd47_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l964_c11_9b1e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_left;
     BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output := BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l973_c21_010e] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_left;
     BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_return_output := BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l961_c11_353a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_left;
     BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output := BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_2a6c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_2a6c_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_6a03 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_6a03_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_75f2 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_75f2_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l967_l961_l975_l964_DUPLICATE_c598 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l967_l961_l975_l964_DUPLICATE_c598_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l967_c11_eb1a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_left;
     BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_return_output := BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l967_l964_DUPLICATE_60df LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l967_l964_DUPLICATE_60df_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l956_c6_d13e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_left;
     BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output := BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l975_c11_661d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_left;
     BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_return_output := BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_cbea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_cbea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c6_d13e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_fc74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_fc74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l961_c11_353a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_5cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_5cff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l964_c11_9b1e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_805f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_eb1a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l975_c11_661d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l973_c21_010e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_75f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_75f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_75f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_75f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l967_l961_l975_l964_DUPLICATE_c598_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l967_l961_l975_l964_DUPLICATE_c598_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l967_l961_l975_l964_DUPLICATE_c598_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l967_l961_l975_l964_DUPLICATE_c598_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_2a6c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_2a6c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_2a6c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_2a6c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_bd47_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_bd47_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_bd47_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l961_l975_l964_l956_DUPLICATE_bd47_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l967_l964_DUPLICATE_60df_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l967_l964_DUPLICATE_60df_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_6a03_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_6a03_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_6a03_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l967_l961_l964_l956_DUPLICATE_6a03_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l970_c30_f07a_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l967_c7_805f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l956_c1_02c9] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l975_c7_df82] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l967_c7_805f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l975_c7_df82] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_return_output;

     -- n8_MUX[uxn_opcodes_h_l967_c7_805f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l967_c7_805f_cond <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_805f_cond;
     n8_MUX_uxn_opcodes_h_l967_c7_805f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_805f_iftrue;
     n8_MUX_uxn_opcodes_h_l967_c7_805f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l967_c7_805f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l967_c7_805f_return_output := n8_MUX_uxn_opcodes_h_l967_c7_805f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l975_c7_df82] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l967_c7_805f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_return_output := result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_return_output;

     -- t8_MUX[uxn_opcodes_h_l964_c7_5cff] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l964_c7_5cff_cond <= VAR_t8_MUX_uxn_opcodes_h_l964_c7_5cff_cond;
     t8_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue;
     t8_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output := t8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l957_c3_0a25_uxn_opcodes_h_l957_c3_0a25_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l956_c1_02c9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse := VAR_n8_MUX_uxn_opcodes_h_l967_c7_805f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l975_c7_df82_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l975_c7_df82_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l975_c7_df82_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l967_c7_805f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l967_c7_805f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse := VAR_t8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l964_c7_5cff] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_cond;
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_return_output := result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;

     -- n8_MUX[uxn_opcodes_h_l964_c7_5cff] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l964_c7_5cff_cond <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_5cff_cond;
     n8_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue;
     n8_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output := n8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;

     -- printf_uxn_opcodes_h_l957_c3_0a25[uxn_opcodes_h_l957_c3_0a25] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l957_c3_0a25_uxn_opcodes_h_l957_c3_0a25_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l957_c3_0a25_uxn_opcodes_h_l957_c3_0a25_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l964_c7_5cff] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l967_c7_805f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l964_c7_5cff] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l967_c7_805f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_return_output;

     -- t8_MUX[uxn_opcodes_h_l961_c7_fc74] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l961_c7_fc74_cond <= VAR_t8_MUX_uxn_opcodes_h_l961_c7_fc74_cond;
     t8_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue;
     t8_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output := t8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l967_c7_805f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse := VAR_n8_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_805f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_805f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_805f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse := VAR_t8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l961_c7_fc74] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l961_c7_fc74] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_cond;
     result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_return_output := result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l964_c7_5cff] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l964_c7_5cff] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l961_c7_fc74] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;

     -- n8_MUX[uxn_opcodes_h_l961_c7_fc74] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l961_c7_fc74_cond <= VAR_n8_MUX_uxn_opcodes_h_l961_c7_fc74_cond;
     n8_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue;
     n8_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output := n8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;

     -- t8_MUX[uxn_opcodes_h_l956_c2_cbea] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l956_c2_cbea_cond <= VAR_t8_MUX_uxn_opcodes_h_l956_c2_cbea_cond;
     t8_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue;
     t8_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output := t8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l964_c7_5cff] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse := VAR_n8_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l964_c7_5cff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l961_c7_fc74] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l956_c2_cbea] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l961_c7_fc74] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l956_c2_cbea] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_cond;
     result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_return_output := result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_return_output;

     -- n8_MUX[uxn_opcodes_h_l956_c2_cbea] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l956_c2_cbea_cond <= VAR_n8_MUX_uxn_opcodes_h_l956_c2_cbea_cond;
     n8_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue;
     n8_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output := n8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l956_c2_cbea] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l961_c7_fc74] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l956_c2_cbea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l961_c7_fc74_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l956_c2_cbea] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l956_c2_cbea] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l956_c2_cbea] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l952_l981_DUPLICATE_8b0f LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l952_l981_DUPLICATE_8b0f_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4e73(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c2_cbea_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c2_cbea_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c2_cbea_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c2_cbea_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c2_cbea_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l952_l981_DUPLICATE_8b0f_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l952_l981_DUPLICATE_8b0f_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
