-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity ovr_0CLK_61914e8d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ovr_0CLK_61914e8d;
architecture arch of ovr_0CLK_61914e8d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l302_c6_b64a]
signal BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l302_c2_559a]
signal n8_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l302_c2_559a]
signal t8_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l302_c2_559a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l302_c2_559a]
signal result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l302_c2_559a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l302_c2_559a]
signal result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l302_c2_559a]
signal result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l302_c2_559a]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l302_c2_559a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l302_c2_559a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l302_c2_559a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l315_c11_1f9c]
signal BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l315_c7_7eb5]
signal n8_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l315_c7_7eb5]
signal t8_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l315_c7_7eb5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l315_c7_7eb5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l315_c7_7eb5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l315_c7_7eb5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l315_c7_7eb5]
signal result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l318_c11_e510]
signal BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l318_c7_73c7]
signal n8_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l318_c7_73c7]
signal t8_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l318_c7_73c7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l318_c7_73c7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l318_c7_73c7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l318_c7_73c7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l318_c7_73c7]
signal result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l320_c30_5599]
signal sp_relative_shift_uxn_opcodes_h_l320_c30_5599_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l320_c30_5599_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l320_c30_5599_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l320_c30_5599_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l325_c11_e824]
signal BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l325_c7_4f43]
signal n8_MUX_uxn_opcodes_h_l325_c7_4f43_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l325_c7_4f43_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l325_c7_4f43]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l325_c7_4f43]
signal result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l325_c7_4f43]
signal result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l325_c7_4f43]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l331_c11_0e6a]
signal BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l331_c7_6c61]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l331_c7_6c61]
signal result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l331_c7_6c61]
signal result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e848( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a
BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_left,
BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_right,
BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output);

-- n8_MUX_uxn_opcodes_h_l302_c2_559a
n8_MUX_uxn_opcodes_h_l302_c2_559a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l302_c2_559a_cond,
n8_MUX_uxn_opcodes_h_l302_c2_559a_iftrue,
n8_MUX_uxn_opcodes_h_l302_c2_559a_iffalse,
n8_MUX_uxn_opcodes_h_l302_c2_559a_return_output);

-- t8_MUX_uxn_opcodes_h_l302_c2_559a
t8_MUX_uxn_opcodes_h_l302_c2_559a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l302_c2_559a_cond,
t8_MUX_uxn_opcodes_h_l302_c2_559a_iftrue,
t8_MUX_uxn_opcodes_h_l302_c2_559a_iffalse,
t8_MUX_uxn_opcodes_h_l302_c2_559a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a
result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a
result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a
result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a
result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a
result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_cond,
result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a
result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a
result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c
BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_left,
BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_right,
BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_return_output);

-- n8_MUX_uxn_opcodes_h_l315_c7_7eb5
n8_MUX_uxn_opcodes_h_l315_c7_7eb5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l315_c7_7eb5_cond,
n8_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue,
n8_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse,
n8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output);

-- t8_MUX_uxn_opcodes_h_l315_c7_7eb5
t8_MUX_uxn_opcodes_h_l315_c7_7eb5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l315_c7_7eb5_cond,
t8_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue,
t8_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse,
t8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5
result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5
result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5
result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5
result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_cond,
result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510
BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_left,
BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_right,
BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_return_output);

-- n8_MUX_uxn_opcodes_h_l318_c7_73c7
n8_MUX_uxn_opcodes_h_l318_c7_73c7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l318_c7_73c7_cond,
n8_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue,
n8_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse,
n8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output);

-- t8_MUX_uxn_opcodes_h_l318_c7_73c7
t8_MUX_uxn_opcodes_h_l318_c7_73c7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l318_c7_73c7_cond,
t8_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue,
t8_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse,
t8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7
result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7
result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7
result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7
result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_cond,
result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_return_output);

-- sp_relative_shift_uxn_opcodes_h_l320_c30_5599
sp_relative_shift_uxn_opcodes_h_l320_c30_5599 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l320_c30_5599_ins,
sp_relative_shift_uxn_opcodes_h_l320_c30_5599_x,
sp_relative_shift_uxn_opcodes_h_l320_c30_5599_y,
sp_relative_shift_uxn_opcodes_h_l320_c30_5599_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824
BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_left,
BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_right,
BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_return_output);

-- n8_MUX_uxn_opcodes_h_l325_c7_4f43
n8_MUX_uxn_opcodes_h_l325_c7_4f43 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l325_c7_4f43_cond,
n8_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue,
n8_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse,
n8_MUX_uxn_opcodes_h_l325_c7_4f43_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43
result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43
result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_cond,
result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43
result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a
BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_left,
BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_right,
BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61
result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61
result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_cond,
result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output,
 n8_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
 t8_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_return_output,
 n8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output,
 t8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_return_output,
 n8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output,
 t8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_return_output,
 sp_relative_shift_uxn_opcodes_h_l320_c30_5599_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_return_output,
 n8_MUX_uxn_opcodes_h_l325_c7_4f43_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l307_c3_ab79 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l312_c3_0672 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l316_c3_0fd5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l325_c7_4f43_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l322_c3_1918 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l320_c30_5599_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l320_c30_5599_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l320_c30_5599_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l320_c30_5599_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l325_c7_4f43_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l328_c3_7fab : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l326_c3_2aed : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l332_c3_888f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l331_c7_6c61_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l302_l315_l331_DUPLICATE_a744_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l318_l315_DUPLICATE_97ea_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l325_l315_DUPLICATE_ff56_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l318_l325_l315_l331_DUPLICATE_1ffa_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l337_l298_DUPLICATE_5915_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l307_c3_ab79 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l307_c3_ab79;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_right := to_unsigned(3, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l316_c3_0fd5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l316_c3_0fd5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l332_c3_888f := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l332_c3_888f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l312_c3_0672 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l312_c3_0672;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l320_c30_5599_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_right := to_unsigned(4, 3);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l326_c3_2aed := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l326_c3_2aed;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l328_c3_7fab := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l328_c3_7fab;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l322_c3_1918 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l322_c3_1918;
     VAR_sp_relative_shift_uxn_opcodes_h_l320_c30_5599_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l320_c30_5599_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l302_c2_559a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse := n8;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l302_c2_559a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l325_c11_e824] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_left;
     BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_return_output := BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l331_c7_6c61] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l331_c7_6c61_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l320_c30_5599] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l320_c30_5599_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l320_c30_5599_ins;
     sp_relative_shift_uxn_opcodes_h_l320_c30_5599_x <= VAR_sp_relative_shift_uxn_opcodes_h_l320_c30_5599_x;
     sp_relative_shift_uxn_opcodes_h_l320_c30_5599_y <= VAR_sp_relative_shift_uxn_opcodes_h_l320_c30_5599_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l320_c30_5599_return_output := sp_relative_shift_uxn_opcodes_h_l320_c30_5599_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l302_c6_b64a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_left;
     BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output := BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l331_c11_0e6a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_left;
     BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_return_output := BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l302_c2_559a_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l318_l315_DUPLICATE_97ea LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l318_l315_DUPLICATE_97ea_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l302_l315_l331_DUPLICATE_a744 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l302_l315_l331_DUPLICATE_a744_return_output := result.u8_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l302_c2_559a_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l318_l325_l315_l331_DUPLICATE_1ffa LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l318_l325_l315_l331_DUPLICATE_1ffa_return_output := result.is_opc_done;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l302_c2_559a_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l315_c11_1f9c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_left;
     BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_return_output := BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l318_c11_e510] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_left;
     BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_return_output := BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l302_c2_559a_return_output := result.is_pc_updated;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l325_l315_DUPLICATE_ff56 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l325_l315_DUPLICATE_ff56_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l302_c2_559a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l302_c2_559a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l302_c6_b64a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l315_c7_7eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l315_c7_7eb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_1f9c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l318_c7_73c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l318_c7_73c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l318_c11_e510_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l325_c7_4f43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_e824_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l331_c11_0e6a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l325_l315_DUPLICATE_ff56_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l325_l315_DUPLICATE_ff56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l318_l325_l315_l331_DUPLICATE_1ffa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l318_l325_l315_l331_DUPLICATE_1ffa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l318_l325_l315_l331_DUPLICATE_1ffa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l318_l325_l315_l331_DUPLICATE_1ffa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l318_l315_DUPLICATE_97ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l318_l315_DUPLICATE_97ea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l302_l315_l331_DUPLICATE_a744_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l302_l315_l331_DUPLICATE_a744_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l302_l315_l331_DUPLICATE_a744_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l302_c2_559a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l302_c2_559a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l302_c2_559a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l302_c2_559a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l331_c7_6c61_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l320_c30_5599_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l318_c7_73c7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l325_c7_4f43] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output;

     -- t8_MUX[uxn_opcodes_h_l318_c7_73c7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l318_c7_73c7_cond <= VAR_t8_MUX_uxn_opcodes_h_l318_c7_73c7_cond;
     t8_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue;
     t8_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output := t8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_return_output;

     -- n8_MUX[uxn_opcodes_h_l325_c7_4f43] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l325_c7_4f43_cond <= VAR_n8_MUX_uxn_opcodes_h_l325_c7_4f43_cond;
     n8_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue;
     n8_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l325_c7_4f43_return_output := n8_MUX_uxn_opcodes_h_l325_c7_4f43_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l331_c7_6c61] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l331_c7_6c61] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_cond;
     result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_return_output := result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l331_c7_6c61] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse := VAR_n8_MUX_uxn_opcodes_h_l325_c7_4f43_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l331_c7_6c61_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l325_c7_4f43_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l331_c7_6c61_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l331_c7_6c61_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse := VAR_t8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l315_c7_7eb5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l325_c7_4f43] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_cond;
     result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_return_output := result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_return_output;

     -- t8_MUX[uxn_opcodes_h_l315_c7_7eb5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l315_c7_7eb5_cond <= VAR_t8_MUX_uxn_opcodes_h_l315_c7_7eb5_cond;
     t8_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue;
     t8_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output := t8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l325_c7_4f43] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l325_c7_4f43] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l318_c7_73c7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;

     -- n8_MUX[uxn_opcodes_h_l318_c7_73c7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l318_c7_73c7_cond <= VAR_n8_MUX_uxn_opcodes_h_l318_c7_73c7_cond;
     n8_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue;
     n8_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output := n8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_4f43_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l325_c7_4f43_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l325_c7_4f43_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l302_c2_559a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l318_c7_73c7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l315_c7_7eb5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;

     -- t8_MUX[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l302_c2_559a_cond <= VAR_t8_MUX_uxn_opcodes_h_l302_c2_559a_cond;
     t8_MUX_uxn_opcodes_h_l302_c2_559a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l302_c2_559a_iftrue;
     t8_MUX_uxn_opcodes_h_l302_c2_559a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l302_c2_559a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l302_c2_559a_return_output := t8_MUX_uxn_opcodes_h_l302_c2_559a_return_output;

     -- n8_MUX[uxn_opcodes_h_l315_c7_7eb5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l315_c7_7eb5_cond <= VAR_n8_MUX_uxn_opcodes_h_l315_c7_7eb5_cond;
     n8_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue;
     n8_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output := n8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l318_c7_73c7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l318_c7_73c7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_return_output := result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l302_c2_559a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l318_c7_73c7_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l302_c2_559a_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l315_c7_7eb5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;

     -- n8_MUX[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l302_c2_559a_cond <= VAR_n8_MUX_uxn_opcodes_h_l302_c2_559a_cond;
     n8_MUX_uxn_opcodes_h_l302_c2_559a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l302_c2_559a_iftrue;
     n8_MUX_uxn_opcodes_h_l302_c2_559a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l302_c2_559a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l302_c2_559a_return_output := n8_MUX_uxn_opcodes_h_l302_c2_559a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l315_c7_7eb5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output := result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l315_c7_7eb5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l302_c2_559a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_7eb5_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_return_output := result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l302_c2_559a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l337_l298_DUPLICATE_5915 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l337_l298_DUPLICATE_5915_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e848(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l302_c2_559a_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l302_c2_559a_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l337_l298_DUPLICATE_5915_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l337_l298_DUPLICATE_5915_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
