-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sft_0CLK_46cced44 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sft_0CLK_46cced44;
architecture arch of sft_0CLK_46cced44 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2213_c6_1473]
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2213_c2_1914]
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2213_c2_1914]
signal n8_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2213_c2_1914]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2213_c2_1914]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2213_c2_1914]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2213_c2_1914]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2213_c2_1914]
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2213_c2_1914]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2213_c2_1914]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2213_c2_1914]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2213_c2_1914]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2213_c2_1914]
signal t8_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2226_c11_0962]
signal BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2226_c7_1be6]
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2226_c7_1be6]
signal n8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2226_c7_1be6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2226_c7_1be6]
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2226_c7_1be6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2226_c7_1be6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2226_c7_1be6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2226_c7_1be6]
signal t8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2229_c11_bd07]
signal BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2229_c7_f0a3]
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2229_c7_f0a3]
signal n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2229_c7_f0a3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2229_c7_f0a3]
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2229_c7_f0a3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2229_c7_f0a3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2229_c7_f0a3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2229_c7_f0a3]
signal t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2231_c30_6f78]
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2233_c11_4347]
signal BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2233_c7_bffa]
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2233_c7_bffa]
signal n8_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2233_c7_bffa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2233_c7_bffa]
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2233_c7_bffa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2233_c7_bffa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2233_c7_bffa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : unsigned(3 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2236_c18_9209]
signal BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_return_output : unsigned(7 downto 0);

-- BIN_OP_SR[uxn_opcodes_h_l2236_c11_7215]
signal BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_left : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_right : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_return_output : unsigned(7 downto 0);

-- CONST_SR_4[uxn_opcodes_h_l2236_c34_32f7]
signal CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7_x : unsigned(7 downto 0);
signal CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7_return_output : unsigned(7 downto 0);

-- BIN_OP_SL[uxn_opcodes_h_l2236_c11_e1ae]
signal BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_left : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_right : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_opc_done := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_left,
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_right,
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2213_c2_1914
tmp8_MUX_uxn_opcodes_h_l2213_c2_1914 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_cond,
tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue,
tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse,
tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output);

-- n8_MUX_uxn_opcodes_h_l2213_c2_1914
n8_MUX_uxn_opcodes_h_l2213_c2_1914 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2213_c2_1914_cond,
n8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue,
n8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse,
n8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_cond,
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_return_output);

-- t8_MUX_uxn_opcodes_h_l2213_c2_1914
t8_MUX_uxn_opcodes_h_l2213_c2_1914 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2213_c2_1914_cond,
t8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue,
t8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse,
t8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_left,
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_right,
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6
tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond,
tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue,
tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse,
tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output);

-- n8_MUX_uxn_opcodes_h_l2226_c7_1be6
n8_MUX_uxn_opcodes_h_l2226_c7_1be6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond,
n8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue,
n8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse,
n8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output);

-- t8_MUX_uxn_opcodes_h_l2226_c7_1be6
t8_MUX_uxn_opcodes_h_l2226_c7_1be6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond,
t8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue,
t8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse,
t8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_left,
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_right,
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3
tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond,
tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue,
tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse,
tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output);

-- n8_MUX_uxn_opcodes_h_l2229_c7_f0a3
n8_MUX_uxn_opcodes_h_l2229_c7_f0a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond,
n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue,
n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse,
n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output);

-- t8_MUX_uxn_opcodes_h_l2229_c7_f0a3
t8_MUX_uxn_opcodes_h_l2229_c7_f0a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond,
t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue,
t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse,
t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78
sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_ins,
sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_x,
sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_y,
sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_left,
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_right,
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa
tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_cond,
tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue,
tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse,
tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output);

-- n8_MUX_uxn_opcodes_h_l2233_c7_bffa
n8_MUX_uxn_opcodes_h_l2233_c7_bffa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2233_c7_bffa_cond,
n8_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue,
n8_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse,
n8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_cond,
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209
BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_left,
BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_right,
BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_return_output);

-- BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215
BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215 : entity work.BIN_OP_SR_uint8_t_uint8_t_0CLK_25d197a7 port map (
BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_left,
BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_right,
BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_return_output);

-- CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7
CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7 : entity work.CONST_SR_4_uint8_t_0CLK_de264c78 port map (
CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7_x,
CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7_return_output);

-- BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae
BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae : entity work.BIN_OP_SL_uint8_t_uint8_t_0CLK_10d8c973 port map (
BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_left,
BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_right,
BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output,
 tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
 n8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
 t8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output,
 tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output,
 n8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output,
 t8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output,
 tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output,
 n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output,
 t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output,
 sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_return_output,
 tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output,
 n8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_return_output,
 BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_return_output,
 CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7_return_output,
 BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2218_c3_0c7f : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_1404 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_1914_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2227_c3_f26e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_6de1 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2238_c3_fa27 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_left : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_right : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7_x : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_ebd1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_0756_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2226_l2233_DUPLICATE_2bc2_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_cda1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_c895_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2243_l2209_DUPLICATE_677d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2218_c3_0c7f := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2218_c3_0c7f;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_1404 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_1404;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_right := to_unsigned(15, 8);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_6de1 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_6de1;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2238_c3_fa27 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2238_c3_fa27;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2227_c3_f26e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2227_c3_f26e;
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_left := VAR_phase;
     VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_left := t8;
     VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7_x := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse := tmp8;
     -- BIN_OP_AND[uxn_opcodes_h_l2236_c18_9209] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_left;
     BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_return_output := BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_0756 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_0756_return_output := result.is_stack_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2213_c2_1914_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_c895 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_c895_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2213_c2_1914_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2229_c11_bd07] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_left;
     BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output := BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2213_c6_1473] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_left;
     BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output := BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2226_l2233_DUPLICATE_2bc2 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2226_l2233_DUPLICATE_2bc2_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l2231_c30_6f78] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_ins;
     sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_x;
     sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_return_output := sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2233_c11_4347] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_left;
     BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_return_output := BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2213_c2_1914_return_output := result.is_pc_updated;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2213_c2_1914_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_ebd1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_ebd1_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_cda1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_cda1_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2226_c11_0962] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_left;
     BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output := BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output;

     -- CONST_SR_4[uxn_opcodes_h_l2236_c34_32f7] LATENCY=0
     -- Inputs
     CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7_x <= VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7_x;
     -- Outputs
     VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7_return_output := CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7_return_output;

     -- Submodule level 1
     VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_right := VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_9209_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_1914_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_1914_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_1473_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_0962_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_bd07_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_bffa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_4347_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2226_l2233_DUPLICATE_2bc2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2226_l2233_DUPLICATE_2bc2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_cda1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_cda1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_cda1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_0756_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_0756_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2226_l2229_l2233_DUPLICATE_0756_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_c895_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_c895_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_ebd1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_ebd1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_ebd1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2226_l2229_l2213_l2233_DUPLICATE_ebd1_return_output;
     VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_right := VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_32f7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2213_c2_1914_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2213_c2_1914_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2213_c2_1914_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2213_c2_1914_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_6f78_return_output;
     -- t8_MUX[uxn_opcodes_h_l2229_c7_f0a3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond <= VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond;
     t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue;
     t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output := t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2233_c7_bffa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2233_c7_bffa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2233_c7_bffa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;

     -- BIN_OP_SR[uxn_opcodes_h_l2236_c11_7215] LATENCY=0
     -- Inputs
     BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_left <= VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_left;
     BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_right <= VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_right;
     -- Outputs
     VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_return_output := BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_return_output;

     -- n8_MUX[uxn_opcodes_h_l2233_c7_bffa] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2233_c7_bffa_cond <= VAR_n8_MUX_uxn_opcodes_h_l2233_c7_bffa_cond;
     n8_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue;
     n8_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output := n8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2233_c7_bffa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;

     -- Submodule level 2
     VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_left := VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_7215_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2229_c7_f0a3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2229_c7_f0a3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;

     -- BIN_OP_SL[uxn_opcodes_h_l2236_c11_e1ae] LATENCY=0
     -- Inputs
     BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_left <= VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_left;
     BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_right <= VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_right;
     -- Outputs
     VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_return_output := BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_return_output;

     -- t8_MUX[uxn_opcodes_h_l2226_c7_1be6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond <= VAR_t8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond;
     t8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue;
     t8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output := t8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;

     -- n8_MUX[uxn_opcodes_h_l2229_c7_f0a3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond <= VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond;
     n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue;
     n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output := n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2229_c7_f0a3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2229_c7_f0a3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_e1ae_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;
     -- t8_MUX[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2213_c2_1914_cond <= VAR_t8_MUX_uxn_opcodes_h_l2213_c2_1914_cond;
     t8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue;
     t8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output := t8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2233_c7_bffa] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output := result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;

     -- n8_MUX[uxn_opcodes_h_l2226_c7_1be6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond <= VAR_n8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond;
     n8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue;
     n8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output := n8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2226_c7_1be6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2226_c7_1be6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2233_c7_bffa] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_cond;
     tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output := tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2226_c7_1be6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2226_c7_1be6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_bffa_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2229_c7_f0a3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;

     -- n8_MUX[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2213_c2_1914_cond <= VAR_n8_MUX_uxn_opcodes_h_l2213_c2_1914_cond;
     n8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue;
     n8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output := n8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2229_c7_f0a3] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_cond;
     tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output := tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_f0a3_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2226_c7_1be6] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_cond;
     tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output := tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2226_c7_1be6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_1be6_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_cond;
     tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output := tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2213_c2_1914] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_return_output := result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;

     -- Submodule level 7
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_1914_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2243_l2209_DUPLICATE_677d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2243_l2209_DUPLICATE_677d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_1914_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_1914_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2243_l2209_DUPLICATE_677d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2243_l2209_DUPLICATE_677d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
