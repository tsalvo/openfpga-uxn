-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity rot_0CLK_b288bfb7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end rot_0CLK_b288bfb7;
architecture arch of rot_0CLK_b288bfb7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2640_c6_62b0]
signal BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2640_c2_0664]
signal l8_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2640_c2_0664]
signal t8_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2640_c2_0664]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2640_c2_0664]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2640_c2_0664]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2640_c2_0664]
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2640_c2_0664]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2640_c2_0664]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2640_c2_0664]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2640_c2_0664]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2640_c2_0664]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2640_c2_0664]
signal n8_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2653_c11_dfb1]
signal BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2653_c7_b77a]
signal l8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2653_c7_b77a]
signal t8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2653_c7_b77a]
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2653_c7_b77a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2653_c7_b77a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2653_c7_b77a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2653_c7_b77a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2653_c7_b77a]
signal n8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2656_c11_0ce6]
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2656_c7_a9e8]
signal l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2656_c7_a9e8]
signal t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2656_c7_a9e8]
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2656_c7_a9e8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2656_c7_a9e8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2656_c7_a9e8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2656_c7_a9e8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2656_c7_a9e8]
signal n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2660_c11_9f4d]
signal BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2660_c7_76fc]
signal l8_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2660_c7_76fc]
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2660_c7_76fc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2660_c7_76fc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2660_c7_76fc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2660_c7_76fc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2660_c7_76fc]
signal n8_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2662_c30_432e]
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2667_c11_5b3e]
signal BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2667_c7_4b47]
signal l8_MUX_uxn_opcodes_h_l2667_c7_4b47_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2667_c7_4b47]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2667_c7_4b47]
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2667_c7_4b47]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2667_c7_4b47]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2673_c11_afa4]
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2673_c7_5bf1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2673_c7_5bf1]
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2673_c7_5bf1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output : unsigned(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_375c( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_vram_write := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.sp_relative_shift := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_left,
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_right,
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output);

-- l8_MUX_uxn_opcodes_h_l2640_c2_0664
l8_MUX_uxn_opcodes_h_l2640_c2_0664 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2640_c2_0664_cond,
l8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue,
l8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse,
l8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output);

-- t8_MUX_uxn_opcodes_h_l2640_c2_0664
t8_MUX_uxn_opcodes_h_l2640_c2_0664 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2640_c2_0664_cond,
t8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue,
t8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse,
t8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_cond,
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_return_output);

-- n8_MUX_uxn_opcodes_h_l2640_c2_0664
n8_MUX_uxn_opcodes_h_l2640_c2_0664 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2640_c2_0664_cond,
n8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue,
n8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse,
n8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_left,
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_right,
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output);

-- l8_MUX_uxn_opcodes_h_l2653_c7_b77a
l8_MUX_uxn_opcodes_h_l2653_c7_b77a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond,
l8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue,
l8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse,
l8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output);

-- t8_MUX_uxn_opcodes_h_l2653_c7_b77a
t8_MUX_uxn_opcodes_h_l2653_c7_b77a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond,
t8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue,
t8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse,
t8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output);

-- n8_MUX_uxn_opcodes_h_l2653_c7_b77a
n8_MUX_uxn_opcodes_h_l2653_c7_b77a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond,
n8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue,
n8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse,
n8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_left,
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_right,
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output);

-- l8_MUX_uxn_opcodes_h_l2656_c7_a9e8
l8_MUX_uxn_opcodes_h_l2656_c7_a9e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond,
l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue,
l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse,
l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output);

-- t8_MUX_uxn_opcodes_h_l2656_c7_a9e8
t8_MUX_uxn_opcodes_h_l2656_c7_a9e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond,
t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue,
t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse,
t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output);

-- n8_MUX_uxn_opcodes_h_l2656_c7_a9e8
n8_MUX_uxn_opcodes_h_l2656_c7_a9e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond,
n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue,
n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse,
n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_left,
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_right,
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_return_output);

-- l8_MUX_uxn_opcodes_h_l2660_c7_76fc
l8_MUX_uxn_opcodes_h_l2660_c7_76fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2660_c7_76fc_cond,
l8_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue,
l8_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse,
l8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_cond,
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output);

-- n8_MUX_uxn_opcodes_h_l2660_c7_76fc
n8_MUX_uxn_opcodes_h_l2660_c7_76fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2660_c7_76fc_cond,
n8_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue,
n8_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse,
n8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2662_c30_432e
sp_relative_shift_uxn_opcodes_h_l2662_c30_432e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_ins,
sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_x,
sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_y,
sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_left,
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_right,
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_return_output);

-- l8_MUX_uxn_opcodes_h_l2667_c7_4b47
l8_MUX_uxn_opcodes_h_l2667_c7_4b47 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2667_c7_4b47_cond,
l8_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue,
l8_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse,
l8_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_cond,
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_left,
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_right,
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 l8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output,
 l8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
 t8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
 n8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output,
 l8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output,
 t8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output,
 n8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output,
 l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output,
 t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output,
 n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_return_output,
 l8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output,
 n8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output,
 sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_return_output,
 l8_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2650_c3_48f7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2645_c3_e0d1 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_0664_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2654_c3_791e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2657_c3_d15c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2664_c3_b10c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_76fc_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_4b47_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_9fee : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2669_c3_a205 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_a572 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2673_c7_5bf1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_2695_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2667_l2660_l2656_l2653_DUPLICATE_b9be_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_34c8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_e98f_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_375c_uxn_opcodes_h_l2679_l2636_DUPLICATE_b708_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_a572 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_a572;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2650_c3_48f7 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2650_c3_48f7;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_right := to_unsigned(3, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2669_c3_a205 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2669_c3_a205;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2657_c3_d15c := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2657_c3_d15c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_9fee := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_9fee;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2654_c3_791e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2654_c3_791e;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2664_c3_b10c := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2664_c3_b10c;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2645_c3_e0d1 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2645_c3_e0d1;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_ins := VAR_ins;
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse := l8;
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_left := VAR_phase;
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2656_c11_0ce6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2640_c2_0664_return_output := result.is_vram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2640_c2_0664_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2660_c11_9f4d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2640_c6_62b0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_34c8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_34c8_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2667_c11_5b3e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_e98f LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_e98f_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l2662_c30_432e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_ins;
     sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_x;
     sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_return_output := sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_2695 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_2695_return_output := result.u8_value;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2640_c2_0664_return_output := result.is_pc_updated;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2640_c2_0664_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2673_c11_afa4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2667_l2660_l2656_l2653_DUPLICATE_b9be LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2667_l2660_l2656_l2653_DUPLICATE_b9be_return_output := result.is_opc_done;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2673_c7_5bf1] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2673_c7_5bf1_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2653_c11_dfb1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_left;
     BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output := BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output;

     -- Submodule level 1
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_0664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_0664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_0664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_62b0_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_dfb1_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0ce6_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_76fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_76fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_9f4d_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_4b47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_5b3e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_afa4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_e98f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_e98f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_e98f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2667_l2660_l2656_l2653_DUPLICATE_b9be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2667_l2660_l2656_l2653_DUPLICATE_b9be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2667_l2660_l2656_l2653_DUPLICATE_b9be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2667_l2660_l2656_l2653_DUPLICATE_b9be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2667_l2660_l2656_l2653_DUPLICATE_b9be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_34c8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_34c8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_34c8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_2695_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_2695_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_2695_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_2695_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2640_c2_0664_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2640_c2_0664_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2640_c2_0664_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2640_c2_0664_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2673_c7_5bf1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_432e_return_output;
     -- t8_MUX[uxn_opcodes_h_l2656_c7_a9e8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond <= VAR_t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond;
     t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue;
     t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output := t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2673_c7_5bf1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output := result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2660_c7_76fc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2667_c7_4b47] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2673_c7_5bf1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;

     -- l8_MUX[uxn_opcodes_h_l2667_c7_4b47] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2667_c7_4b47_cond <= VAR_l8_MUX_uxn_opcodes_h_l2667_c7_4b47_cond;
     l8_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue;
     l8_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output := l8_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;

     -- n8_MUX[uxn_opcodes_h_l2660_c7_76fc] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2660_c7_76fc_cond <= VAR_n8_MUX_uxn_opcodes_h_l2660_c7_76fc_cond;
     n8_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue;
     n8_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output := n8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2673_c7_5bf1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;

     -- Submodule level 2
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_5bf1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;
     -- l8_MUX[uxn_opcodes_h_l2660_c7_76fc] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2660_c7_76fc_cond <= VAR_l8_MUX_uxn_opcodes_h_l2660_c7_76fc_cond;
     l8_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue;
     l8_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output := l8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;

     -- t8_MUX[uxn_opcodes_h_l2653_c7_b77a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond <= VAR_t8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond;
     t8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue;
     t8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output := t8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;

     -- n8_MUX[uxn_opcodes_h_l2656_c7_a9e8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond;
     n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue;
     n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output := n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2667_c7_4b47] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output := result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2667_c7_4b47] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2660_c7_76fc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2667_c7_4b47] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2656_c7_a9e8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;

     -- Submodule level 3
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_4b47_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;
     -- n8_MUX[uxn_opcodes_h_l2653_c7_b77a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond <= VAR_n8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond;
     n8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue;
     n8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output := n8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2660_c7_76fc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2660_c7_76fc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;

     -- t8_MUX[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2640_c2_0664_cond <= VAR_t8_MUX_uxn_opcodes_h_l2640_c2_0664_cond;
     t8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue;
     t8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output := t8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;

     -- l8_MUX[uxn_opcodes_h_l2656_c7_a9e8] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond <= VAR_l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond;
     l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue;
     l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output := l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2656_c7_a9e8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2653_c7_b77a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2660_c7_76fc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output := result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;

     -- Submodule level 4
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_76fc_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2656_c7_a9e8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2653_c7_b77a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;

     -- l8_MUX[uxn_opcodes_h_l2653_c7_b77a] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond <= VAR_l8_MUX_uxn_opcodes_h_l2653_c7_b77a_cond;
     l8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue;
     l8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output := l8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2656_c7_a9e8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2656_c7_a9e8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;

     -- n8_MUX[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2640_c2_0664_cond <= VAR_n8_MUX_uxn_opcodes_h_l2640_c2_0664_cond;
     n8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue;
     n8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output := n8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;

     -- Submodule level 5
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_a9e8_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2653_c7_b77a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2653_c7_b77a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2653_c7_b77a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;

     -- l8_MUX[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2640_c2_0664_cond <= VAR_l8_MUX_uxn_opcodes_h_l2640_c2_0664_cond;
     l8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue;
     l8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output := l8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;

     -- Submodule level 6
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_b77a_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_return_output := result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2640_c2_0664] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_375c_uxn_opcodes_h_l2679_l2636_DUPLICATE_b708 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_375c_uxn_opcodes_h_l2679_l2636_DUPLICATE_b708_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_375c(
     result,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_0664_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_0664_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_375c_uxn_opcodes_h_l2679_l2636_DUPLICATE_b708_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_375c_uxn_opcodes_h_l2679_l2636_DUPLICATE_b708_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
