-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 17
entity VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_0CLK_83e31706 is
port(
 elem_val : in unsigned(7 downto 0);
 ref_toks_0 : in uint8_t_8;
 var_dim_0 : in unsigned(2 downto 0);
 return_output : out uint8_t_array_8_t);
end VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_0CLK_83e31706;
architecture arch of VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_0CLK_83e31706 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_return_output : unsigned(0 downto 0);

-- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe]
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_cond : unsigned(0 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_iftrue : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_iffalse : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_return_output : unsigned(0 downto 0);

-- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1]
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_cond : unsigned(0 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_iftrue : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_iffalse : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_return_output : unsigned(0 downto 0);

-- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736]
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_cond : unsigned(0 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_iftrue : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_iffalse : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_return_output : unsigned(0 downto 0);

-- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7]
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_cond : unsigned(0 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_iftrue : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_iffalse : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_return_output : unsigned(0 downto 0);

-- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d]
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_cond : unsigned(0 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_iftrue : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_iffalse : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_return_output : unsigned(0 downto 0);

-- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96]
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_cond : unsigned(0 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_iftrue : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_iffalse : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_return_output : unsigned(0 downto 0);

-- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410]
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_cond : unsigned(0 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_iftrue : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_iffalse : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_left : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_return_output : unsigned(0 downto 0);

-- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495]
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_cond : unsigned(0 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_iftrue : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_iffalse : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_return_output : unsigned(7 downto 0);

function CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_ab7c( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return uint8_t_array_8_t is
 
  variable base : uint8_t_array_8_t; 
  variable return_output : uint8_t_array_8_t;
begin
      base.data(2) := ref_toks_0;
      base.data(5) := ref_toks_1;
      base.data(1) := ref_toks_2;
      base.data(4) := ref_toks_3;
      base.data(7) := ref_toks_4;
      base.data(3) := ref_toks_5;
      base.data(0) := ref_toks_6;
      base.data(6) := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e : entity work.BIN_OP_EQ_uint3_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_return_output);

-- rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_cond,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_iftrue,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_iffalse,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08 : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_return_output);

-- rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_cond,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_iftrue,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_iffalse,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c : entity work.BIN_OP_EQ_uint3_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_return_output);

-- rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_cond,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_iftrue,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_iffalse,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_return_output);

-- rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_cond,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_iftrue,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_iffalse,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_return_output);

-- rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_cond,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_iftrue,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_iffalse,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0 : entity work.BIN_OP_EQ_uint3_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_return_output);

-- rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_cond,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_iftrue,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_iffalse,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c : entity work.BIN_OP_EQ_uint3_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_return_output);

-- rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_cond,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_iftrue,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_iffalse,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5 : entity work.BIN_OP_EQ_uint3_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_return_output);

-- rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_cond,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_iftrue,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_iffalse,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 elem_val,
 ref_toks_0,
 var_dim_0,
 -- All submodule outputs
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_return_output,
 rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_return_output,
 rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_return_output,
 rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_return_output,
 rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_return_output,
 rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_return_output,
 rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_return_output,
 rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_return_output,
 rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_elem_val : unsigned(7 downto 0);
 variable VAR_ref_toks_0 : uint8_t_8;
 variable VAR_var_dim_0 : unsigned(2 downto 0);
 variable VAR_return_output : uint8_t_array_8_t;
 variable VAR_base : uint8_t_8;
 variable VAR_rv : uint8_t_array_8_t;
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_9fc4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_e259_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_29c3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_c72e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_787f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_4294_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_bb59_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_b0cc_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_left : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_ab7c_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_795e_return_output : uint8_t_array_8_t;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_right := to_unsigned(6, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_elem_val := elem_val;
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_iftrue := VAR_elem_val;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_iftrue := VAR_elem_val;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_iftrue := VAR_elem_val;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_iftrue := VAR_elem_val;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_iftrue := VAR_elem_val;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_iftrue := VAR_elem_val;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_iftrue := VAR_elem_val;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_iftrue := VAR_elem_val;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_left := VAR_var_dim_0;
     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_2_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_9fc4] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_9fc4_return_output := VAR_ref_toks_0(2);

     -- CONST_REF_RD_uint8_t_uint8_t_8_7_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_787f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_787f_return_output := VAR_ref_toks_0(7);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_5_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_e259] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_e259_return_output := VAR_ref_toks_0(5);

     -- CONST_REF_RD_uint8_t_uint8_t_8_3_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_4294] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_4294_return_output := VAR_ref_toks_0(3);

     -- CONST_REF_RD_uint8_t_uint8_t_8_4_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_c72e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_c72e_return_output := VAR_ref_toks_0(4);

     -- CONST_REF_RD_uint8_t_uint8_t_8_0_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_bb59] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_bb59_return_output := VAR_ref_toks_0(0);

     -- CONST_REF_RD_uint8_t_uint8_t_8_1_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_29c3] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_29c3_return_output := VAR_ref_toks_0(1);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_8_6_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_b0cc] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_b0cc_return_output := VAR_ref_toks_0(6);

     -- Submodule level 1
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l25_c5_a09e_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l31_c5_8f08_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l37_c5_d67c_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l43_c5_5b8d_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l49_c5_768d_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l55_c5_02b0_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l61_c5_a16c_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l67_c5_76c5_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l21_c15_bb59_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l17_c15_29c3_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l15_c15_9fc4_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l20_c15_4294_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l18_c15_c72e_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l16_c15_e259_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l22_c15_b0cc_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_8_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l19_c15_787f_return_output;
     -- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7] LATENCY=0
     -- Inputs
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_cond <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_cond;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_iftrue <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_iftrue;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_iffalse <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_iffalse;
     -- Outputs
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_return_output := rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_return_output;

     -- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410] LATENCY=0
     -- Inputs
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_cond <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_cond;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_iftrue <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_iftrue;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_iffalse <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_iffalse;
     -- Outputs
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_return_output := rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_return_output;

     -- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96] LATENCY=0
     -- Inputs
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_cond <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_cond;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_iftrue <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_iftrue;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_iffalse <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_iffalse;
     -- Outputs
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_return_output := rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_return_output;

     -- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe] LATENCY=0
     -- Inputs
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_cond <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_cond;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_iftrue <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_iftrue;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_iffalse <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_iffalse;
     -- Outputs
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_return_output := rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_return_output;

     -- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d] LATENCY=0
     -- Inputs
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_cond <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_cond;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_iftrue <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_iftrue;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_iffalse <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_iffalse;
     -- Outputs
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_return_output := rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_return_output;

     -- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736] LATENCY=0
     -- Inputs
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_cond <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_cond;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_iftrue <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_iftrue;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_iffalse <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_iffalse;
     -- Outputs
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_return_output := rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_return_output;

     -- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1] LATENCY=0
     -- Inputs
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_cond <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_cond;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_iftrue <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_iftrue;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_iffalse <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_iffalse;
     -- Outputs
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_return_output := rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_return_output;

     -- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495] LATENCY=0
     -- Inputs
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_cond <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_cond;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_iftrue <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_iftrue;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_iffalse <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_iffalse;
     -- Outputs
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_return_output := rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_return_output;

     -- Submodule level 2
     -- CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_ab7c[VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_795e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_ab7c_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_795e_return_output := CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_ab7c(
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l24_c2_46fe_return_output,
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l30_c2_74b1_return_output,
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l36_c2_d736_return_output,
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l42_c2_b6b7_return_output,
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l48_c2_566d_return_output,
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l54_c2_aa96_return_output,
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l60_c2_0410_return_output,
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l66_c2_c495_return_output);

     -- Submodule level 3
     VAR_return_output := VAR_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_ab7c_VAR_REF_ASSIGN_uint8_t_uint8_t_8_VAR_52b8_c_l73_c10_795e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
