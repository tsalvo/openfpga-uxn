-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 48
entity ldr_0CLK_f74745d5 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr_0CLK_f74745d5;
architecture arch of ldr_0CLK_f74745d5 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1600_c6_081f]
signal BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1600_c2_9ec7]
signal t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1600_c2_9ec7]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1600_c2_9ec7]
signal result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1600_c2_9ec7]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1600_c2_9ec7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1600_c2_9ec7]
signal result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1600_c2_9ec7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1600_c2_9ec7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1600_c2_9ec7]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1600_c2_9ec7]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1600_c2_9ec7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1600_c2_9ec7]
signal tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1613_c11_0935]
signal BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1613_c7_d773]
signal t8_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1613_c7_d773]
signal result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1613_c7_d773]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1613_c7_d773]
signal result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1613_c7_d773]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1613_c7_d773]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1613_c7_d773]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1613_c7_d773]
signal tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1616_c11_c395]
signal BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1616_c7_0c68]
signal t8_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1616_c7_0c68]
signal result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1616_c7_0c68]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1616_c7_0c68]
signal result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1616_c7_0c68]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1616_c7_0c68]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1616_c7_0c68]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1616_c7_0c68]
signal tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1618_c30_ef39]
signal sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1619_c22_24b1]
signal BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1621_c11_7fbb]
signal BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1621_c7_e699]
signal result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1621_c7_e699]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1621_c7_e699]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1621_c7_e699]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1621_c7_e699]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1621_c7_e699]
signal tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1624_c11_7020]
signal BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1624_c7_2642]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1624_c7_2642]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1624_c7_2642]
signal result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1624_c7_2642]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_return_output : unsigned(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1624_c7_2642]
signal tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_return_output : unsigned(7 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_d9be( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_vram_write := ref_toks_1;
      base.u16_value := ref_toks_2;
      base.is_pc_updated := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_index_flipped := ref_toks_9;
      base.sp_relative_shift := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f
BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_left,
BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_right,
BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output);

-- t8_MUX_uxn_opcodes_h_l1600_c2_9ec7
t8_MUX_uxn_opcodes_h_l1600_c2_9ec7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond,
t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue,
t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse,
t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7
result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7
result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond,
result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7
result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7
result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7
result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond,
result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7
result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7
result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7
result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7
tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond,
tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue,
tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse,
tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935
BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_left,
BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_right,
BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output);

-- t8_MUX_uxn_opcodes_h_l1613_c7_d773
t8_MUX_uxn_opcodes_h_l1613_c7_d773 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1613_c7_d773_cond,
t8_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue,
t8_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse,
t8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773
result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_cond,
result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773
result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773
result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_cond,
result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773
result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773
result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1613_c7_d773
tmp8_MUX_uxn_opcodes_h_l1613_c7_d773 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_cond,
tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue,
tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse,
tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395
BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_left,
BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_right,
BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output);

-- t8_MUX_uxn_opcodes_h_l1616_c7_0c68
t8_MUX_uxn_opcodes_h_l1616_c7_0c68 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1616_c7_0c68_cond,
t8_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue,
t8_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse,
t8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68
result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_cond,
result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68
result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68
result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_cond,
result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68
result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68
result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68
tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_cond,
tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue,
tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse,
tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39
sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_ins,
sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_x,
sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_y,
sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1
BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_left,
BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_right,
BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb
BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_left,
BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_right,
BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699
result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_cond,
result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699
result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699
result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699
result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1621_c7_e699
tmp8_MUX_uxn_opcodes_h_l1621_c7_e699 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_cond,
tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue,
tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse,
tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020
BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_left,
BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_right,
BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642
result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642
result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642
result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_cond,
result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1624_c7_2642
tmp8_MUX_uxn_opcodes_h_l1624_c7_2642 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_cond,
tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue,
tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse,
tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output,
 t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
 tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output,
 t8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_return_output,
 tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output,
 t8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output,
 tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output,
 sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_return_output,
 tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_return_output,
 tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1610_c3_45b0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1605_c3_6d27 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1614_c3_5769 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1619_c3_8758 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1619_c27_0232_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1622_c3_a664 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1627_c3_676b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1613_l1616_l1600_DUPLICATE_fac7_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1616_l1613_l1600_l1624_l1621_DUPLICATE_c030_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_38d5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_172b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1613_l1621_DUPLICATE_2ad1_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1624_l1616_l1621_DUPLICATE_38c5_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d9be_uxn_opcodes_h_l1632_l1596_DUPLICATE_a32a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1627_c3_676b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1627_c3_676b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1605_c3_6d27 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1605_c3_6d27;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1614_c3_5769 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1614_c3_5769;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1622_c3_a664 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1622_c3_a664;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1610_c3_45b0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1610_c3_45b0;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1600_c6_081f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1600_c2_9ec7_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_172b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_172b_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1613_c11_0935] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_left;
     BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output := BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1613_l1616_l1600_DUPLICATE_fac7 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1613_l1616_l1600_DUPLICATE_fac7_return_output := result.u16_value;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1616_l1613_l1600_l1624_l1621_DUPLICATE_c030 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1616_l1613_l1600_l1624_l1621_DUPLICATE_c030_return_output := result.u8_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1624_l1616_l1621_DUPLICATE_38c5 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1624_l1616_l1621_DUPLICATE_38c5_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1613_l1621_DUPLICATE_2ad1 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1613_l1621_DUPLICATE_2ad1_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1624_c11_7020] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_left;
     BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_return_output := BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1600_c2_9ec7_return_output := result.is_stack_index_flipped;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1600_c2_9ec7_return_output := result.is_ram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1600_c2_9ec7_return_output := result.is_pc_updated;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1619_c27_0232] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1619_c27_0232_return_output := CAST_TO_int8_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1616_c11_c395] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_left;
     BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output := BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1621_c11_7fbb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_left;
     BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_return_output := BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_38d5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_38d5_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l1618_c30_ef39] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_ins;
     sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_x;
     sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_return_output := sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1600_c6_081f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1613_c7_d773_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1613_c11_0935_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1616_c7_0c68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1616_c11_c395_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1621_c11_7fbb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1624_c11_7020_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1619_c27_0232_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1613_l1621_DUPLICATE_2ad1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1613_l1621_DUPLICATE_2ad1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1613_l1616_l1600_DUPLICATE_fac7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1613_l1616_l1600_DUPLICATE_fac7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1613_l1616_l1600_DUPLICATE_fac7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_38d5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_38d5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_38d5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_38d5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_172b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_172b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_172b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1613_l1624_l1616_l1621_DUPLICATE_172b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1624_l1616_l1621_DUPLICATE_38c5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1624_l1616_l1621_DUPLICATE_38c5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1624_l1616_l1621_DUPLICATE_38c5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1616_l1613_l1600_l1624_l1621_DUPLICATE_c030_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1616_l1613_l1600_l1624_l1621_DUPLICATE_c030_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1616_l1613_l1600_l1624_l1621_DUPLICATE_c030_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1616_l1613_l1600_l1624_l1621_DUPLICATE_c030_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1616_l1613_l1600_l1624_l1621_DUPLICATE_c030_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1600_c2_9ec7_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1600_c2_9ec7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1600_c2_9ec7_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1600_c2_9ec7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_ef39_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l1624_c7_2642] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_cond;
     tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_return_output := tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1624_c7_2642] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_return_output := result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1619_c22_24b1] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_return_output;

     -- t8_MUX[uxn_opcodes_h_l1616_c7_0c68] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1616_c7_0c68_cond <= VAR_t8_MUX_uxn_opcodes_h_l1616_c7_0c68_cond;
     t8_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue;
     t8_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output := t8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1621_c7_e699] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1624_c7_2642] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1624_c7_2642] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1624_c7_2642] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1619_c3_8758 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1619_c22_24b1_return_output)),16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1624_c7_2642_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1624_c7_2642_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1621_c7_e699_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1624_c7_2642_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1624_c7_2642_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1624_c7_2642_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1619_c3_8758;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1621_c7_e699] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1621_c7_e699] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_cond;
     tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_return_output := tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1616_c7_0c68] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;

     -- t8_MUX[uxn_opcodes_h_l1613_c7_d773] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1613_c7_d773_cond <= VAR_t8_MUX_uxn_opcodes_h_l1613_c7_d773_cond;
     t8_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue;
     t8_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output := t8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1621_c7_e699] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1616_c7_0c68] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output := result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1621_c7_e699] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1621_c7_e699] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_return_output := result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1621_c7_e699_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1621_c7_e699_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1621_c7_e699_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1621_c7_e699_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1621_c7_e699_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1613_c7_d773] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1616_c7_0c68] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output := result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1616_c7_0c68] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1616_c7_0c68] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;

     -- t8_MUX[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond <= VAR_t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond;
     t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue;
     t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output := t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1616_c7_0c68] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1613_c7_d773] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output := result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1616_c7_0c68] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_cond;
     tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output := tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1616_c7_0c68_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1613_c7_d773] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1613_c7_d773] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_cond;
     tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output := tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1613_c7_d773] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1613_c7_d773] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output := result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output := result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1613_c7_d773] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1613_c7_d773_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output := result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond;
     tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output := tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1600_c2_9ec7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;

     -- Submodule level 6
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_d9be_uxn_opcodes_h_l1632_l1596_DUPLICATE_a32a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d9be_uxn_opcodes_h_l1632_l1596_DUPLICATE_a32a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_d9be(
     result,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1600_c2_9ec7_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d9be_uxn_opcodes_h_l1632_l1596_DUPLICATE_a32a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d9be_uxn_opcodes_h_l1632_l1596_DUPLICATE_a32a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
