-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 61
entity ldr2_0CLK_b7cf2331 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr2_0CLK_b7cf2331;
architecture arch of ldr2_0CLK_b7cf2331 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8_high : unsigned(7 downto 0);
signal REG_COMB_tmp8_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1638_c6_523a]
signal BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1638_c2_30fc]
signal result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1638_c2_30fc]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1638_c2_30fc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1638_c2_30fc]
signal result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(15 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1638_c2_30fc]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1638_c2_30fc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1638_c2_30fc]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1638_c2_30fc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1638_c2_30fc]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1638_c2_30fc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1638_c2_30fc]
signal t8_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(7 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l1638_c2_30fc]
signal tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l1638_c2_30fc]
signal tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1651_c11_9436]
signal BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1651_c7_0aa2]
signal result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1651_c7_0aa2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1651_c7_0aa2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : signed(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1651_c7_0aa2]
signal result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1651_c7_0aa2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1651_c7_0aa2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1651_c7_0aa2]
signal t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(7 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l1651_c7_0aa2]
signal tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l1651_c7_0aa2]
signal tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1652_c30_ce1a]
signal sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1654_c11_f7e2]
signal BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1654_c7_4c1c]
signal result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1654_c7_4c1c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1654_c7_4c1c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : signed(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1654_c7_4c1c]
signal result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1654_c7_4c1c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1654_c7_4c1c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1654_c7_4c1c]
signal t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(7 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l1654_c7_4c1c]
signal tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l1654_c7_4c1c]
signal tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1657_c22_1b91]
signal BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1659_c11_7992]
signal BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1659_c7_13b7]
signal result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1659_c7_13b7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1659_c7_13b7]
signal result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1659_c7_13b7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1659_c7_13b7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l1659_c7_13b7]
signal tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l1659_c7_13b7]
signal tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1660_c22_b6e1]
signal BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_return_output : signed(17 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1660_c22_1cc0]
signal BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_left : signed(17 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_right : signed(1 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_return_output : signed(18 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1662_c11_4672]
signal BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1662_c7_23df]
signal result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1662_c7_23df]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1662_c7_23df]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1662_c7_23df]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l1662_c7_23df]
signal tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l1662_c7_23df]
signal tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1668_c11_3fc8]
signal BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1668_c7_d204]
signal result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1668_c7_d204]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1668_c7_d204]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_return_output : unsigned(0 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l1668_c7_d204]
signal tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_return_output : unsigned(7 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_e482( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.u16_value := ref_toks_4;
      base.is_vram_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_opc_done := ref_toks_8;
      base.is_ram_write := ref_toks_9;
      base.is_stack_write := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a
BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_left,
BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_right,
BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc
result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_cond,
result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc
result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_cond,
result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc
result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc
result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc
result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

-- t8_MUX_uxn_opcodes_h_l1638_c2_30fc
t8_MUX_uxn_opcodes_h_l1638_c2_30fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1638_c2_30fc_cond,
t8_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue,
t8_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse,
t8_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc
tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_cond,
tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc
tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_cond,
tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436
BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_left,
BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_right,
BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2
result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2
result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond,
result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2
result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2
result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output);

-- t8_MUX_uxn_opcodes_h_l1651_c7_0aa2
t8_MUX_uxn_opcodes_h_l1651_c7_0aa2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond,
t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue,
t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse,
t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2
tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond,
tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2
tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond,
tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a
sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_ins,
sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_x,
sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_y,
sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2
BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_left,
BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_right,
BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c
result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c
result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond,
result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c
result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c
result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output);

-- t8_MUX_uxn_opcodes_h_l1654_c7_4c1c
t8_MUX_uxn_opcodes_h_l1654_c7_4c1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond,
t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue,
t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse,
t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c
tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond,
tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c
tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond,
tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91
BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_left,
BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_right,
BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992
BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_left,
BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_right,
BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7
result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_cond,
result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7
result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_cond,
result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7
result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7
result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7
tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_cond,
tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7
tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_cond,
tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1
BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_left,
BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_right,
BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0
BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0 : entity work.BIN_OP_PLUS_int18_t_int2_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_left,
BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_right,
BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672
BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_left,
BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_right,
BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df
result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_cond,
result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df
result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df
result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df
tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_cond,
tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df
tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_cond,
tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8
BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_left,
BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_right,
BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204
result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_cond,
result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204
result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204
tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_cond,
tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8_high,
 tmp8_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
 t8_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output,
 t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output,
 sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output,
 t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1648_c3_2044 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1643_c3_2d0a : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1656_c3_f2b8 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1654_c7_4c1c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1657_c3_49af : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1657_c27_c62e_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1660_c3_c51b : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1660_c27_a1dc_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_left : signed(17 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_right : signed(1 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_return_output : signed(18 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1665_c3_cdad : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_cond : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1670_c3_50fa : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1654_l1651_l1638_l1668_l1659_DUPLICATE_0ce4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1638_l1659_l1651_DUPLICATE_5186_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1654_l1668_l1659_l1651_DUPLICATE_35d8_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1654_l1651_l1668_l1662_l1659_DUPLICATE_bb92_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1654_l1659_l1651_l1662_DUPLICATE_f25b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e482_uxn_opcodes_h_l1675_l1634_DUPLICATE_de5f_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8_high : unsigned(7 downto 0);
variable REG_VAR_tmp8_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8_high := tmp8_high;
  REG_VAR_tmp8_low := tmp8_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1656_c3_f2b8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1656_c3_f2b8;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1643_c3_2d0a := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1643_c3_2d0a;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1670_c3_50fa := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1670_c3_50fa;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1648_c3_2044 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1648_c3_2044;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_right := signed(std_logic_vector(resize(to_unsigned(1, 1), 2)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1665_c3_cdad := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1665_c3_cdad;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue := VAR_previous_ram_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue := VAR_previous_ram_read;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue := VAR_previous_ram_read;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse := t8;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse := tmp8_high;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse := tmp8_low;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1654_l1651_l1668_l1662_l1659_DUPLICATE_bb92 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1654_l1651_l1668_l1662_l1659_DUPLICATE_bb92_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1651_c11_9436] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_left;
     BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output := BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1668_c11_3fc8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1654_c11_f7e2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1638_c2_30fc_return_output := result.is_ram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1638_c2_30fc_return_output := result.is_pc_updated;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1657_c27_c62e] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1657_c27_c62e_return_output := CAST_TO_int8_t_uint8_t(
     VAR_previous_stack_read);

     -- sp_relative_shift[uxn_opcodes_h_l1652_c30_ce1a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_ins;
     sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_x;
     sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_return_output := sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1638_l1659_l1651_DUPLICATE_5186 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1638_l1659_l1651_DUPLICATE_5186_return_output := result.u16_value;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l1654_c7_4c1c] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1654_c7_4c1c_return_output := result.sp_relative_shift;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1638_c2_30fc_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1662_c11_4672] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_left;
     BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_return_output := BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1638_c6_523a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1654_l1659_l1651_l1662_DUPLICATE_f25b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1654_l1659_l1651_l1662_DUPLICATE_f25b_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1654_l1651_l1638_l1668_l1659_DUPLICATE_0ce4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1654_l1651_l1638_l1668_l1659_DUPLICATE_0ce4_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1659_c11_7992] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_left;
     BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_return_output := BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1638_c2_30fc_return_output := result.is_vram_write;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1660_c27_a1dc] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1660_c27_a1dc_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1654_l1668_l1659_l1651_DUPLICATE_35d8 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1654_l1668_l1659_l1651_DUPLICATE_35d8_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1638_c2_30fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1638_c6_523a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1651_c11_9436_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1654_c11_f7e2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1659_c11_7992_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1662_c11_4672_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1668_c11_3fc8_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1657_c27_c62e_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1660_c27_a1dc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1638_l1659_l1651_DUPLICATE_5186_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1638_l1659_l1651_DUPLICATE_5186_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1638_l1659_l1651_DUPLICATE_5186_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1654_l1651_l1668_l1662_l1659_DUPLICATE_bb92_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1654_l1651_l1668_l1662_l1659_DUPLICATE_bb92_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1654_l1651_l1668_l1662_l1659_DUPLICATE_bb92_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1654_l1651_l1668_l1662_l1659_DUPLICATE_bb92_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1654_l1651_l1668_l1662_l1659_DUPLICATE_bb92_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1654_l1659_l1651_l1662_DUPLICATE_f25b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1654_l1659_l1651_l1662_DUPLICATE_f25b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1654_l1659_l1651_l1662_DUPLICATE_f25b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1654_l1659_l1651_l1662_DUPLICATE_f25b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1654_l1668_l1659_l1651_DUPLICATE_35d8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1654_l1668_l1659_l1651_DUPLICATE_35d8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1654_l1668_l1659_l1651_DUPLICATE_35d8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1654_l1668_l1659_l1651_DUPLICATE_35d8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1654_l1651_l1638_l1668_l1659_DUPLICATE_0ce4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1654_l1651_l1638_l1668_l1659_DUPLICATE_0ce4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1654_l1651_l1638_l1668_l1659_DUPLICATE_0ce4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1654_l1651_l1638_l1668_l1659_DUPLICATE_0ce4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1654_l1651_l1638_l1668_l1659_DUPLICATE_0ce4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1638_c2_30fc_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1638_c2_30fc_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1638_c2_30fc_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1638_c2_30fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1654_c7_4c1c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1652_c30_ce1a_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l1668_c7_d204] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_cond;
     tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_return_output := tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1668_c7_d204] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1654_c7_4c1c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1654_c7_4c1c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond <= VAR_t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond;
     t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue;
     t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output := t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1668_c7_d204] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_return_output := result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1657_c22_1b91] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1662_c7_23df] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1660_c22_b6e1] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l1662_c7_23df] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_cond;
     tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_return_output := tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1668_c7_d204] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1657_c3_49af := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1657_c22_1b91_return_output)),16);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_left := VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_b6e1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1668_c7_d204_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1662_c7_23df_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1668_c7_d204_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1668_c7_d204_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l1662_c7_23df_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l1668_c7_d204_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1657_c3_49af;
     -- result_u8_value_MUX[uxn_opcodes_h_l1662_c7_23df] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_return_output := result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_return_output;

     -- t8_MUX[uxn_opcodes_h_l1651_c7_0aa2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond <= VAR_t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond;
     t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue;
     t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output := t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l1662_c7_23df] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_cond;
     tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_return_output := tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1659_c7_13b7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l1659_c7_13b7] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_cond;
     tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output := tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1651_c7_0aa2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1662_c7_23df] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1662_c7_23df] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1660_c22_1cc0] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_return_output;

     -- Submodule level 3
     VAR_result_u16_value_uxn_opcodes_h_l1660_c3_c51b := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1660_c22_1cc0_return_output)),16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1662_c7_23df_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1662_c7_23df_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1662_c7_23df_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l1662_c7_23df_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1660_c3_c51b;
     -- tmp8_low_MUX[uxn_opcodes_h_l1659_c7_13b7] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_cond;
     tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output := tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1659_c7_13b7] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output := result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1654_c7_4c1c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1659_c7_13b7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l1654_c7_4c1c] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond;
     tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output := tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1638_c2_30fc_cond <= VAR_t8_MUX_uxn_opcodes_h_l1638_c2_30fc_cond;
     t8_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue;
     t8_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output := t8_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1659_c7_13b7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output := result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1659_c7_13b7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l1659_c7_13b7_return_output;
     -- tmp8_high_MUX[uxn_opcodes_h_l1651_c7_0aa2] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond;
     tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output := tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1654_c7_4c1c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l1654_c7_4c1c] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond;
     tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output := tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1651_c7_0aa2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1654_c7_4c1c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output := result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1654_c7_4c1c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1654_c7_4c1c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l1654_c7_4c1c_return_output;
     -- tmp8_low_MUX[uxn_opcodes_h_l1651_c7_0aa2] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond;
     tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output := tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_cond;
     tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output := tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1651_c7_0aa2] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output := result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1651_c7_0aa2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1651_c7_0aa2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1651_c7_0aa2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;
     REG_VAR_tmp8_high := VAR_tmp8_high_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l1651_c7_0aa2_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output := result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output := result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l1638_c2_30fc] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_cond;
     tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output := tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;

     -- Submodule level 7
     REG_VAR_tmp8_low := VAR_tmp8_low_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e482_uxn_opcodes_h_l1675_l1634_DUPLICATE_de5f LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e482_uxn_opcodes_h_l1675_l1634_DUPLICATE_de5f_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e482(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1638_c2_30fc_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e482_uxn_opcodes_h_l1675_l1634_DUPLICATE_de5f_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e482_uxn_opcodes_h_l1675_l1634_DUPLICATE_de5f_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8_high <= REG_VAR_tmp8_high;
REG_COMB_tmp8_low <= REG_VAR_tmp8_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8_high <= REG_COMB_tmp8_high;
     tmp8_low <= REG_COMB_tmp8_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
