-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity sub_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub_0CLK_f62d646e;
architecture arch of sub_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2622_c6_1cab]
signal BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2622_c1_898c]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2622_c2_e23d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2622_c2_e23d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2622_c2_e23d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2622_c2_e23d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2622_c2_e23d]
signal result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2622_c2_e23d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2622_c2_e23d]
signal t8_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2622_c2_e23d]
signal n8_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2623_c3_d8b4[uxn_opcodes_h_l2623_c3_d8b4]
signal printf_uxn_opcodes_h_l2623_c3_d8b4_uxn_opcodes_h_l2623_c3_d8b4_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2627_c11_5c93]
signal BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2627_c7_41c8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2627_c7_41c8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2627_c7_41c8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2627_c7_41c8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2627_c7_41c8]
signal result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2627_c7_41c8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2627_c7_41c8]
signal t8_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2627_c7_41c8]
signal n8_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2630_c11_fe09]
signal BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2630_c7_d935]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2630_c7_d935]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2630_c7_d935]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2630_c7_d935]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2630_c7_d935]
signal result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2630_c7_d935]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2630_c7_d935]
signal t8_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2630_c7_d935]
signal n8_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2634_c11_0ee9]
signal BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2634_c7_2568]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2634_c7_2568]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2634_c7_2568]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2634_c7_2568]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2634_c7_2568]
signal result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2634_c7_2568]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2634_c7_2568]
signal n8_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2637_c11_e542]
signal BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2637_c7_f434]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2637_c7_f434]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2637_c7_f434]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2637_c7_f434]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2637_c7_f434]
signal result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2637_c7_f434]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2637_c7_f434]
signal n8_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2640_c30_7b02]
signal sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_return_output : signed(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2643_c21_5bd6]
signal BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2645_c11_b0b7]
signal BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2645_c7_8466]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2645_c7_8466]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2645_c7_8466]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_641b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab
BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_left,
BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_right,
BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d
result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d
result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d
result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d
result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output);

-- t8_MUX_uxn_opcodes_h_l2622_c2_e23d
t8_MUX_uxn_opcodes_h_l2622_c2_e23d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2622_c2_e23d_cond,
t8_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue,
t8_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse,
t8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output);

-- n8_MUX_uxn_opcodes_h_l2622_c2_e23d
n8_MUX_uxn_opcodes_h_l2622_c2_e23d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2622_c2_e23d_cond,
n8_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue,
n8_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse,
n8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output);

-- printf_uxn_opcodes_h_l2623_c3_d8b4_uxn_opcodes_h_l2623_c3_d8b4
printf_uxn_opcodes_h_l2623_c3_d8b4_uxn_opcodes_h_l2623_c3_d8b4 : entity work.printf_uxn_opcodes_h_l2623_c3_d8b4_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2623_c3_d8b4_uxn_opcodes_h_l2623_c3_d8b4_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93
BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_left,
BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_right,
BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8
result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8
result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8
result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8
result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output);

-- t8_MUX_uxn_opcodes_h_l2627_c7_41c8
t8_MUX_uxn_opcodes_h_l2627_c7_41c8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2627_c7_41c8_cond,
t8_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue,
t8_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse,
t8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output);

-- n8_MUX_uxn_opcodes_h_l2627_c7_41c8
n8_MUX_uxn_opcodes_h_l2627_c7_41c8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2627_c7_41c8_cond,
n8_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue,
n8_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse,
n8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09
BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_left,
BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_right,
BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935
result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935
result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935
result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935
result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_cond,
result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935
result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output);

-- t8_MUX_uxn_opcodes_h_l2630_c7_d935
t8_MUX_uxn_opcodes_h_l2630_c7_d935 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2630_c7_d935_cond,
t8_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue,
t8_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse,
t8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output);

-- n8_MUX_uxn_opcodes_h_l2630_c7_d935
n8_MUX_uxn_opcodes_h_l2630_c7_d935 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2630_c7_d935_cond,
n8_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue,
n8_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse,
n8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9
BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_left,
BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_right,
BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568
result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568
result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568
result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568
result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_cond,
result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568
result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output);

-- n8_MUX_uxn_opcodes_h_l2634_c7_2568
n8_MUX_uxn_opcodes_h_l2634_c7_2568 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2634_c7_2568_cond,
n8_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue,
n8_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse,
n8_MUX_uxn_opcodes_h_l2634_c7_2568_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542
BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_left,
BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_right,
BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434
result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434
result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434
result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434
result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_cond,
result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434
result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output);

-- n8_MUX_uxn_opcodes_h_l2637_c7_f434
n8_MUX_uxn_opcodes_h_l2637_c7_f434 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2637_c7_f434_cond,
n8_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue,
n8_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse,
n8_MUX_uxn_opcodes_h_l2637_c7_f434_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02
sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_ins,
sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_x,
sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_y,
sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6
BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_left,
BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_right,
BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7
BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_left,
BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_right,
BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466
result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466
result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466
result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output,
 t8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output,
 n8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output,
 t8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output,
 n8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output,
 t8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output,
 n8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output,
 n8_MUX_uxn_opcodes_h_l2634_c7_2568_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output,
 n8_MUX_uxn_opcodes_h_l2637_c7_f434_return_output,
 sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2624_c3_dcaa : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2622_c2_e23d_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2623_c3_d8b4_uxn_opcodes_h_l2623_c3_d8b4_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2628_c3_ed41 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2627_c7_41c8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2632_c3_9d7a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2634_c7_2568_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2630_c7_d935_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2635_c3_6e19 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2637_c7_f434_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2634_c7_2568_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2642_c3_0c19 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2637_c7_f434_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2637_c7_f434_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_722f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_3396_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_82a6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_1120_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2627_l2645_l2637_l2634_l2630_DUPLICATE_ef61_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2651_l2618_DUPLICATE_b958_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2628_c3_ed41 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2628_c3_ed41;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2635_c3_6e19 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2635_c3_6e19;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2632_c3_9d7a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2632_c3_9d7a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2642_c3_0c19 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2642_c3_0c19;
     VAR_sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_right := to_unsigned(4, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2624_c3_dcaa := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2624_c3_dcaa;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_1120 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_1120_return_output := result.sp_relative_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2637_c7_f434] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2637_c7_f434_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2630_c11_fe09] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_left;
     BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output := BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2645_c11_b0b7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_left;
     BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_return_output := BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2627_l2645_l2637_l2634_l2630_DUPLICATE_ef61 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2627_l2645_l2637_l2634_l2630_DUPLICATE_ef61_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l2640_c30_7b02] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_ins;
     sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_x;
     sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_return_output := sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_return_output;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2643_c21_5bd6] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2634_c11_0ee9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2622_c6_1cab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_left;
     BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output := BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_722f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_722f_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_3396 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_3396_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2627_c11_5c93] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_left;
     BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output := BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2637_c11_e542] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_left;
     BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_return_output := BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_82a6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_82a6_return_output := result.u8_value;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2622_c2_e23d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2622_c2_e23d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c6_1cab_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2627_c7_41c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2627_c7_41c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c11_5c93_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2630_c7_d935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2630_c7_d935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2630_c11_fe09_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2634_c7_2568_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2634_c11_0ee9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2637_c7_f434_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_e542_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2645_c11_b0b7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2643_c21_5bd6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_1120_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_1120_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_1120_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_1120_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_1120_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2627_l2645_l2637_l2634_l2630_DUPLICATE_ef61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2627_l2645_l2637_l2634_l2630_DUPLICATE_ef61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2627_l2645_l2637_l2634_l2630_DUPLICATE_ef61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2627_l2645_l2637_l2634_l2630_DUPLICATE_ef61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2627_l2645_l2637_l2634_l2630_DUPLICATE_ef61_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_722f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_722f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_722f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_722f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_722f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_3396_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_3396_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_3396_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_3396_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2627_l2622_l2645_l2634_l2630_DUPLICATE_3396_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_82a6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_82a6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_82a6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_82a6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2627_l2622_l2637_l2634_l2630_DUPLICATE_82a6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2637_c7_f434_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2640_c30_7b02_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2637_c7_f434] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_return_output := result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2637_c7_f434] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2622_c1_898c] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2637_c7_f434] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2637_c7_f434_cond <= VAR_n8_MUX_uxn_opcodes_h_l2637_c7_f434_cond;
     n8_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue;
     n8_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2637_c7_f434_return_output := n8_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2645_c7_8466] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2637_c7_f434] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2645_c7_8466] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2645_c7_8466] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_return_output;

     -- t8_MUX[uxn_opcodes_h_l2630_c7_d935] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2630_c7_d935_cond <= VAR_t8_MUX_uxn_opcodes_h_l2630_c7_d935_cond;
     t8_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue;
     t8_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output := t8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2623_c3_d8b4_uxn_opcodes_h_l2623_c3_d8b4_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2622_c1_898c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2645_c7_8466_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2645_c7_8466_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2645_c7_8466_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2637_c7_f434] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;

     -- printf_uxn_opcodes_h_l2623_c3_d8b4[uxn_opcodes_h_l2623_c3_d8b4] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2623_c3_d8b4_uxn_opcodes_h_l2623_c3_d8b4_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2623_c3_d8b4_uxn_opcodes_h_l2623_c3_d8b4_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2637_c7_f434] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2637_c7_f434] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2634_c7_2568] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_return_output := result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;

     -- t8_MUX[uxn_opcodes_h_l2627_c7_41c8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2627_c7_41c8_cond <= VAR_t8_MUX_uxn_opcodes_h_l2627_c7_41c8_cond;
     t8_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue;
     t8_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output := t8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2634_c7_2568] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2634_c7_2568] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;

     -- n8_MUX[uxn_opcodes_h_l2634_c7_2568] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2634_c7_2568_cond <= VAR_n8_MUX_uxn_opcodes_h_l2634_c7_2568_cond;
     n8_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue;
     n8_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2634_c7_2568_return_output := n8_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_f434_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;
     -- n8_MUX[uxn_opcodes_h_l2630_c7_d935] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2630_c7_d935_cond <= VAR_n8_MUX_uxn_opcodes_h_l2630_c7_d935_cond;
     n8_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue;
     n8_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output := n8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2630_c7_d935] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_return_output := result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;

     -- t8_MUX[uxn_opcodes_h_l2622_c2_e23d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2622_c2_e23d_cond <= VAR_t8_MUX_uxn_opcodes_h_l2622_c2_e23d_cond;
     t8_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue;
     t8_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output := t8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2630_c7_d935] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2634_c7_2568] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2630_c7_d935] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2634_c7_2568] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2634_c7_2568] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2634_c7_2568_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2627_c7_41c8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2627_c7_41c8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;

     -- n8_MUX[uxn_opcodes_h_l2627_c7_41c8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2627_c7_41c8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2627_c7_41c8_cond;
     n8_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue;
     n8_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output := n8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2630_c7_d935] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2630_c7_d935] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2630_c7_d935] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2627_c7_41c8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2630_c7_d935_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2622_c2_e23d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2627_c7_41c8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2622_c2_e23d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2627_c7_41c8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2627_c7_41c8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2622_c2_e23d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output;

     -- n8_MUX[uxn_opcodes_h_l2622_c2_e23d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2622_c2_e23d_cond <= VAR_n8_MUX_uxn_opcodes_h_l2622_c2_e23d_cond;
     n8_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue;
     n8_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output := n8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c7_41c8_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2622_c2_e23d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2622_c2_e23d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2622_c2_e23d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2651_l2618_DUPLICATE_b958 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2651_l2618_DUPLICATE_b958_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_641b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c2_e23d_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2651_l2618_DUPLICATE_b958_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2651_l2618_DUPLICATE_b958_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
