-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sth2_0CLK_55b6500a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth2_0CLK_55b6500a;
architecture arch of sth2_0CLK_55b6500a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2419_c6_3bab]
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2419_c2_5a62]
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2419_c2_5a62]
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2419_c2_5a62]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2419_c2_5a62]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2419_c2_5a62]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2419_c2_5a62]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2419_c2_5a62]
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2419_c2_5a62]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2419_c2_5a62]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2419_c2_5a62]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2419_c2_5a62]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2432_c11_7074]
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2432_c7_71f2]
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2432_c7_71f2]
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2432_c7_71f2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2432_c7_71f2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2432_c7_71f2]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2432_c7_71f2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2432_c7_71f2]
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2432_c7_71f2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2435_c11_3bea]
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2435_c7_0d9b]
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2435_c7_0d9b]
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2435_c7_0d9b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2435_c7_0d9b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2435_c7_0d9b]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2435_c7_0d9b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2435_c7_0d9b]
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2435_c7_0d9b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2437_c30_9a4b]
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2439_c11_23d4]
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2439_c7_de15]
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2439_c7_de15]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2439_c7_de15]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2439_c7_de15]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2439_c7_de15]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2439_c7_de15]
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2439_c7_de15]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2447_c11_eece]
signal BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2447_c7_bbe7]
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2447_c7_bbe7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2447_c7_bbe7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2447_c7_bbe7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output : unsigned(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_opc_done := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_left,
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_right,
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62
t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_cond,
t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue,
t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse,
t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62
t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_cond,
t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue,
t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse,
t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_cond,
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_left,
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_right,
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2
t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_cond,
t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue,
t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse,
t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2
t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_cond,
t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue,
t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse,
t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_left,
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_right,
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b
t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond,
t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue,
t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse,
t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b
t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond,
t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue,
t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse,
t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b
sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_ins,
sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_x,
sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_y,
sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_left,
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_right,
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2439_c7_de15
t16_low_MUX_uxn_opcodes_h_l2439_c7_de15 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_cond,
t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue,
t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse,
t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_cond,
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_left,
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_right,
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond,
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output,
 t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
 t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output,
 t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output,
 t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output,
 t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output,
 t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output,
 sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_return_output,
 t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2424_c3_58af : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_6c91 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_31ba : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2442_c3_c801 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2444_c3_36bb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2448_c3_f771 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2449_c3_2d4b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_bb8f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_441a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_fd33_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_6dba_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_2147_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_595c_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2454_l2415_DUPLICATE_2b92_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2444_c3_36bb := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2444_c3_36bb;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2424_c3_58af := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2424_c3_58af;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_31ba := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_31ba;
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2449_c3_2d4b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2449_c3_2d4b;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_right := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2442_c3_c801 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2442_c3_c801;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2448_c3_f771 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2448_c3_f771;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_6c91 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_6c91;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_right := to_unsigned(2, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_left := VAR_phase;
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse := t16_high;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse := t16_low;
     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2419_c2_5a62_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_fd33 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_fd33_return_output := result.is_stack_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2419_c2_5a62_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_6dba LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_6dba_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2435_c11_3bea] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_left;
     BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output := BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2419_c2_5a62_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2419_c6_3bab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_left;
     BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output := BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_bb8f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_bb8f_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2439_c11_23d4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2432_c11_7074] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_left;
     BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output := BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_441a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_441a_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l2437_c30_9a4b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_ins;
     sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_x;
     sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_return_output := sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2447_c11_eece] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_left;
     BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_return_output := BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_595c LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_595c_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_2147 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_2147_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_3bab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7074_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3bea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_23d4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_eece_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_2147_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_2147_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_441a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_441a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_441a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_441a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_6dba_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_6dba_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_6dba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_fd33_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_fd33_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_fd33_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_595c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_595c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_bb8f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_bb8f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_bb8f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_bb8f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2419_c2_5a62_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2419_c2_5a62_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2419_c2_5a62_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9a4b_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l2435_c7_0d9b] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond;
     t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output := t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2447_c7_bbe7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output := result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2439_c7_de15] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2447_c7_bbe7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2447_c7_bbe7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2447_c7_bbe7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2439_c7_de15] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_cond;
     t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_return_output := t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2439_c7_de15] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_bbe7_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;
     -- t16_low_MUX[uxn_opcodes_h_l2435_c7_0d9b] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond;
     t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output := t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2432_c7_71f2] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_cond;
     t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output := t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2439_c7_de15] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_return_output := result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2439_c7_de15] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2435_c7_0d9b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2439_c7_de15] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2435_c7_0d9b] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2439_c7_de15] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_de15_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2432_c7_71f2] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2432_c7_71f2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2432_c7_71f2] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_cond;
     t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output := t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2435_c7_0d9b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2435_c7_0d9b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2435_c7_0d9b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_cond;
     t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output := t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2435_c7_0d9b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_0d9b_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2432_c7_71f2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2432_c7_71f2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2432_c7_71f2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2432_c7_71f2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_cond;
     t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output := t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_71f2_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2419_c2_5a62] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output := result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2454_l2415_DUPLICATE_2b92 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2454_l2415_DUPLICATE_2b92_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_5a62_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2454_l2415_DUPLICATE_2b92_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2454_l2415_DUPLICATE_2b92_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
