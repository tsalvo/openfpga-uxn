-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 43
entity inc_0CLK_66ba3dc0 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc_0CLK_66ba3dc0;
architecture arch of inc_0CLK_66ba3dc0 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1284_c6_076c]
signal BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1284_c1_5ec8]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1284_c2_e9a7]
signal t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1284_c2_e9a7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1284_c2_e9a7]
signal result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1284_c2_e9a7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1284_c2_e9a7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1284_c2_e9a7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1284_c2_e9a7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1284_c2_e9a7]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l1285_c3_e03a[uxn_opcodes_h_l1285_c3_e03a]
signal printf_uxn_opcodes_h_l1285_c3_e03a_uxn_opcodes_h_l1285_c3_e03a_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1290_c11_ba23]
signal BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1290_c7_4c0f]
signal t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1290_c7_4c0f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1290_c7_4c0f]
signal result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1290_c7_4c0f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1290_c7_4c0f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1290_c7_4c0f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1290_c7_4c0f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1290_c7_4c0f]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1293_c11_d4cf]
signal BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1293_c7_5c1f]
signal t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1293_c7_5c1f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1293_c7_5c1f]
signal result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1293_c7_5c1f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1293_c7_5c1f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1293_c7_5c1f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1293_c7_5c1f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1293_c7_5c1f]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1297_c32_6961]
signal BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1297_c32_332f]
signal BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1297_c32_e3de]
signal MUX_uxn_opcodes_h_l1297_c32_e3de_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1297_c32_e3de_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1297_c32_e3de_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1297_c32_e3de_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1299_c11_9d54]
signal BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1299_c7_038c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1299_c7_038c]
signal result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1299_c7_038c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1299_c7_038c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1299_c7_038c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1303_c24_1fd6]
signal BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1305_c11_7986]
signal BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1305_c7_e71c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1305_c7_e71c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e56b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_sp_shift := ref_toks_1;
      base.stack_value := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_stack_read := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c
BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_left,
BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_right,
BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_return_output);

-- t8_MUX_uxn_opcodes_h_l1284_c2_e9a7
t8_MUX_uxn_opcodes_h_l1284_c2_e9a7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond,
t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue,
t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse,
t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7
result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7
result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond,
result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7
result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7
result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output);

-- printf_uxn_opcodes_h_l1285_c3_e03a_uxn_opcodes_h_l1285_c3_e03a
printf_uxn_opcodes_h_l1285_c3_e03a_uxn_opcodes_h_l1285_c3_e03a : entity work.printf_uxn_opcodes_h_l1285_c3_e03a_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1285_c3_e03a_uxn_opcodes_h_l1285_c3_e03a_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23
BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_left,
BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_right,
BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output);

-- t8_MUX_uxn_opcodes_h_l1290_c7_4c0f
t8_MUX_uxn_opcodes_h_l1290_c7_4c0f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond,
t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue,
t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse,
t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f
result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f
result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond,
result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f
result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f
result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f
result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf
BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_left,
BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_right,
BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output);

-- t8_MUX_uxn_opcodes_h_l1293_c7_5c1f
t8_MUX_uxn_opcodes_h_l1293_c7_5c1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond,
t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue,
t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse,
t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f
result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f
result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond,
result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f
result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f
result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f
result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961
BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_left,
BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_right,
BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f
BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_left,
BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_right,
BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_return_output);

-- MUX_uxn_opcodes_h_l1297_c32_e3de
MUX_uxn_opcodes_h_l1297_c32_e3de : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1297_c32_e3de_cond,
MUX_uxn_opcodes_h_l1297_c32_e3de_iftrue,
MUX_uxn_opcodes_h_l1297_c32_e3de_iffalse,
MUX_uxn_opcodes_h_l1297_c32_e3de_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54
BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_left,
BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_right,
BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c
result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_cond,
result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6
BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_left,
BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_right,
BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986
BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_left,
BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_right,
BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c
result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c
result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_return_output,
 t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output,
 t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output,
 t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_return_output,
 MUX_uxn_opcodes_h_l1297_c32_e3de_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1287_c3_5f21 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1285_c3_e03a_uxn_opcodes_h_l1285_c3_e03a_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1291_c3_bc8f : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1297_c32_e3de_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1297_c32_e3de_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1297_c32_e3de_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1297_c32_e3de_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_uxn_opcodes_h_l1303_c3_e849 : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1302_c3_9128 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_return_output : unsigned(8 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1290_l1284_l1299_DUPLICATE_1a3c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1290_l1293_l1284_l1299_DUPLICATE_f6b3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1290_l1293_l1284_DUPLICATE_1f59_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1284_DUPLICATE_7d85_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1299_DUPLICATE_8254_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1290_l1293_DUPLICATE_46da_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1293_l1299_DUPLICATE_e42b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l1280_l1310_DUPLICATE_c429_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1302_c3_9128 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1302_c3_9128;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1291_c3_bc8f := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1291_c3_bc8f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_right := to_unsigned(2, 2);
     VAR_BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1287_c3_5f21 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1287_c3_5f21;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_right := to_unsigned(3, 2);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_right := to_unsigned(128, 8);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1297_c32_e3de_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_right := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1297_c32_e3de_iffalse := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1290_l1293_DUPLICATE_46da LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1290_l1293_DUPLICATE_46da_return_output := result.is_stack_read;

     -- BIN_OP_EQ[uxn_opcodes_h_l1299_c11_9d54] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_left;
     BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_return_output := BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1293_l1299_DUPLICATE_e42b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1293_l1299_DUPLICATE_e42b_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1284_c6_076c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1284_DUPLICATE_7d85 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1284_DUPLICATE_7d85_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1293_c11_d4cf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_left;
     BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output := BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l1297_c32_6961] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_left;
     BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_return_output := BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1290_c11_ba23] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_left;
     BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output := BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1305_c11_7986] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_left;
     BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_return_output := BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1303_c24_1fd6] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1290_l1293_l1284_DUPLICATE_1f59 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1290_l1293_l1284_DUPLICATE_1f59_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1299_DUPLICATE_8254 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1299_DUPLICATE_8254_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1290_l1284_l1299_DUPLICATE_1a3c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1290_l1284_l1299_DUPLICATE_1a3c_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1290_l1293_l1284_l1299_DUPLICATE_f6b3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1290_l1293_l1284_l1299_DUPLICATE_f6b3_return_output := result.stack_value;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1297_c32_6961_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c6_076c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1290_c11_ba23_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1293_c11_d4cf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1299_c11_9d54_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1305_c11_7986_return_output;
     VAR_result_stack_value_uxn_opcodes_h_l1303_c3_e849 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1303_c24_1fd6_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1290_l1293_l1284_DUPLICATE_1f59_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1290_l1293_l1284_DUPLICATE_1f59_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1290_l1293_l1284_DUPLICATE_1f59_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1299_DUPLICATE_8254_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1299_DUPLICATE_8254_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1299_DUPLICATE_8254_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1299_DUPLICATE_8254_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1290_l1284_l1299_DUPLICATE_1a3c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1290_l1284_l1299_DUPLICATE_1a3c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1290_l1284_l1299_DUPLICATE_1a3c_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1290_l1293_DUPLICATE_46da_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1290_l1293_DUPLICATE_46da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1284_DUPLICATE_7d85_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1284_DUPLICATE_7d85_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1284_DUPLICATE_7d85_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1290_l1305_l1293_l1284_DUPLICATE_7d85_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1293_l1299_DUPLICATE_e42b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1293_l1299_DUPLICATE_e42b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1290_l1293_l1284_l1299_DUPLICATE_f6b3_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1290_l1293_l1284_l1299_DUPLICATE_f6b3_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1290_l1293_l1284_l1299_DUPLICATE_f6b3_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1290_l1293_l1284_l1299_DUPLICATE_f6b3_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue := VAR_result_stack_value_uxn_opcodes_h_l1303_c3_e849;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1305_c7_e71c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1299_c7_038c] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_return_output := result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1297_c32_332f] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_left;
     BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_return_output := BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1284_c1_5ec8] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1293_c7_5c1f] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1299_c7_038c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1299_c7_038c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1305_c7_e71c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1293_c7_5c1f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond;
     t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue;
     t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output := t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1297_c32_e3de_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1297_c32_332f_return_output;
     VAR_printf_uxn_opcodes_h_l1285_c3_e03a_uxn_opcodes_h_l1285_c3_e03a_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1284_c1_5ec8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1299_c7_038c_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1305_c7_e71c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1299_c7_038c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1299_c7_038c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1299_c7_038c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1290_c7_4c0f] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1293_c7_5c1f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;

     -- printf_uxn_opcodes_h_l1285_c3_e03a[uxn_opcodes_h_l1285_c3_e03a] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1285_c3_e03a_uxn_opcodes_h_l1285_c3_e03a_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1285_c3_e03a_uxn_opcodes_h_l1285_c3_e03a_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- MUX[uxn_opcodes_h_l1297_c32_e3de] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1297_c32_e3de_cond <= VAR_MUX_uxn_opcodes_h_l1297_c32_e3de_cond;
     MUX_uxn_opcodes_h_l1297_c32_e3de_iftrue <= VAR_MUX_uxn_opcodes_h_l1297_c32_e3de_iftrue;
     MUX_uxn_opcodes_h_l1297_c32_e3de_iffalse <= VAR_MUX_uxn_opcodes_h_l1297_c32_e3de_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1297_c32_e3de_return_output := MUX_uxn_opcodes_h_l1297_c32_e3de_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1293_c7_5c1f] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output := result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1290_c7_4c0f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond;
     t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue;
     t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output := t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1293_c7_5c1f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1299_c7_038c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue := VAR_MUX_uxn_opcodes_h_l1297_c32_e3de_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1299_c7_038c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1299_c7_038c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;
     -- result_stack_value_MUX[uxn_opcodes_h_l1290_c7_4c0f] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output := result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1293_c7_5c1f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1284_c2_e9a7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond <= VAR_t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond;
     t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue;
     t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output := t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1290_c7_4c0f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1284_c2_e9a7] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1290_c7_4c0f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1293_c7_5c1f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1293_c7_5c1f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1293_c7_5c1f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1284_c2_e9a7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1290_c7_4c0f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1284_c2_e9a7] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output := result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1284_c2_e9a7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1290_c7_4c0f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1290_c7_4c0f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1290_c7_4c0f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1284_c2_e9a7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1284_c2_e9a7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1284_c2_e9a7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l1280_l1310_DUPLICATE_c429 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l1280_l1310_DUPLICATE_c429_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e56b(
     result,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1284_c2_e9a7_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l1280_l1310_DUPLICATE_c429_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l1280_l1310_DUPLICATE_c429_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
