-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 42
entity nip_0CLK_6481cb28 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip_0CLK_6481cb28;
architecture arch of nip_0CLK_6481cb28 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1405_c6_056c]
signal BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1405_c1_246e]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1405_c2_24aa]
signal t8_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1405_c2_24aa]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1405_c2_24aa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1405_c2_24aa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1405_c2_24aa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1405_c2_24aa]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1405_c2_24aa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1405_c2_24aa]
signal result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1406_c3_7745[uxn_opcodes_h_l1406_c3_7745]
signal printf_uxn_opcodes_h_l1406_c3_7745_uxn_opcodes_h_l1406_c3_7745_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1411_c11_a566]
signal BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1411_c7_a63d]
signal t8_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1411_c7_a63d]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1411_c7_a63d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1411_c7_a63d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1411_c7_a63d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1411_c7_a63d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1411_c7_a63d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1411_c7_a63d]
signal result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1414_c11_0eb3]
signal BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1414_c7_1a71]
signal t8_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1414_c7_1a71]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1414_c7_1a71]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1414_c7_1a71]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1414_c7_1a71]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1414_c7_1a71]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1414_c7_1a71]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1414_c7_1a71]
signal result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(7 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1418_c32_7880]
signal BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1418_c32_c41c]
signal BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1418_c32_79e3]
signal MUX_uxn_opcodes_h_l1418_c32_79e3_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1418_c32_79e3_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1418_c32_79e3_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1418_c32_79e3_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1420_c11_e011]
signal BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1420_c7_7f85]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1420_c7_7f85]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1420_c7_7f85]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1420_c7_7f85]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1420_c7_7f85]
signal result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1426_c11_5bf9]
signal BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1426_c7_fc7f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1426_c7_fc7f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_28d7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : signed;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_read := ref_toks_1;
      base.sp_relative_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_sp_shift := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.stack_value := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c
BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_left,
BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_right,
BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_return_output);

-- t8_MUX_uxn_opcodes_h_l1405_c2_24aa
t8_MUX_uxn_opcodes_h_l1405_c2_24aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1405_c2_24aa_cond,
t8_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue,
t8_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse,
t8_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa
result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa
result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa
result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa
result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa
result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa
result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_cond,
result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output);

-- printf_uxn_opcodes_h_l1406_c3_7745_uxn_opcodes_h_l1406_c3_7745
printf_uxn_opcodes_h_l1406_c3_7745_uxn_opcodes_h_l1406_c3_7745 : entity work.printf_uxn_opcodes_h_l1406_c3_7745_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1406_c3_7745_uxn_opcodes_h_l1406_c3_7745_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566
BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_left,
BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_right,
BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output);

-- t8_MUX_uxn_opcodes_h_l1411_c7_a63d
t8_MUX_uxn_opcodes_h_l1411_c7_a63d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1411_c7_a63d_cond,
t8_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue,
t8_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse,
t8_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d
result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d
result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d
result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d
result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d
result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_cond,
result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3
BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_left,
BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_right,
BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output);

-- t8_MUX_uxn_opcodes_h_l1414_c7_1a71
t8_MUX_uxn_opcodes_h_l1414_c7_1a71 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1414_c7_1a71_cond,
t8_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue,
t8_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse,
t8_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71
result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71
result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71
result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71
result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71
result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71
result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_cond,
result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880
BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_left,
BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_right,
BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c
BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_left,
BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_right,
BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_return_output);

-- MUX_uxn_opcodes_h_l1418_c32_79e3
MUX_uxn_opcodes_h_l1418_c32_79e3 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1418_c32_79e3_cond,
MUX_uxn_opcodes_h_l1418_c32_79e3_iftrue,
MUX_uxn_opcodes_h_l1418_c32_79e3_iffalse,
MUX_uxn_opcodes_h_l1418_c32_79e3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011
BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_left,
BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_right,
BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85
result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85
result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85
result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85
result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_cond,
result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9
BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_left,
BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_right,
BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f
result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f
result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_return_output,
 t8_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output,
 t8_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output,
 t8_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_return_output,
 MUX_uxn_opcodes_h_l1418_c32_79e3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1408_c3_104a : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1406_c3_7745_uxn_opcodes_h_l1406_c3_7745_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1412_c3_9a35 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1418_c32_79e3_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1418_c32_79e3_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1418_c32_79e3_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1418_c32_79e3_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1423_c3_ad03 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1414_l1405_l1411_DUPLICATE_4950_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1414_l1405_l1426_l1411_DUPLICATE_4bc8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1405_l1420_l1411_DUPLICATE_4440_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1414_l1405_l1420_l1411_DUPLICATE_6452_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1414_l1411_DUPLICATE_e6de_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1414_l1426_l1420_l1411_DUPLICATE_9565_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1414_l1420_DUPLICATE_5fa0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_28d7_uxn_opcodes_h_l1401_l1431_DUPLICATE_3816_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_right := to_unsigned(1, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_right := to_unsigned(128, 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1418_c32_79e3_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1423_c3_ad03 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1423_c3_ad03;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1412_c3_9a35 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1412_c3_9a35;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_right := to_unsigned(4, 3);
     VAR_MUX_uxn_opcodes_h_l1418_c32_79e3_iffalse := resize(to_signed(-1, 2), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1408_c3_104a := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1408_c3_104a;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_iffalse := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1420_c11_e011] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_left;
     BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_return_output := BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1405_c6_056c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1405_l1420_l1411_DUPLICATE_4440 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1405_l1420_l1411_DUPLICATE_4440_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1414_l1426_l1420_l1411_DUPLICATE_9565 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1414_l1426_l1420_l1411_DUPLICATE_9565_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1414_l1420_DUPLICATE_5fa0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1414_l1420_DUPLICATE_5fa0_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1414_c11_0eb3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1411_c11_a566] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_left;
     BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output := BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1414_l1411_DUPLICATE_e6de LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1414_l1411_DUPLICATE_e6de_return_output := result.is_stack_read;

     -- BIN_OP_EQ[uxn_opcodes_h_l1426_c11_5bf9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1414_l1405_l1420_l1411_DUPLICATE_6452 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1414_l1405_l1420_l1411_DUPLICATE_6452_return_output := result.stack_value;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1414_l1405_l1411_DUPLICATE_4950 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1414_l1405_l1411_DUPLICATE_4950_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1414_l1405_l1426_l1411_DUPLICATE_4bc8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1414_l1405_l1426_l1411_DUPLICATE_4bc8_return_output := result.is_stack_write;

     -- BIN_OP_AND[uxn_opcodes_h_l1418_c32_7880] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_left;
     BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_return_output := BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1418_c32_7880_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1405_c2_24aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1405_c6_056c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1411_c7_a63d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1411_c11_a566_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1414_c7_1a71_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1414_c11_0eb3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1420_c11_e011_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_5bf9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1414_l1405_l1411_DUPLICATE_4950_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1414_l1405_l1411_DUPLICATE_4950_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1414_l1405_l1411_DUPLICATE_4950_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1414_l1426_l1420_l1411_DUPLICATE_9565_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1414_l1426_l1420_l1411_DUPLICATE_9565_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1414_l1426_l1420_l1411_DUPLICATE_9565_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1414_l1426_l1420_l1411_DUPLICATE_9565_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1405_l1420_l1411_DUPLICATE_4440_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1405_l1420_l1411_DUPLICATE_4440_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1405_l1420_l1411_DUPLICATE_4440_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1414_l1411_DUPLICATE_e6de_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1414_l1411_DUPLICATE_e6de_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1414_l1405_l1426_l1411_DUPLICATE_4bc8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1414_l1405_l1426_l1411_DUPLICATE_4bc8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1414_l1405_l1426_l1411_DUPLICATE_4bc8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1414_l1405_l1426_l1411_DUPLICATE_4bc8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1414_l1420_DUPLICATE_5fa0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1414_l1420_DUPLICATE_5fa0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1414_l1405_l1420_l1411_DUPLICATE_6452_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1414_l1405_l1420_l1411_DUPLICATE_6452_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1414_l1405_l1420_l1411_DUPLICATE_6452_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1414_l1405_l1420_l1411_DUPLICATE_6452_return_output;
     -- result_is_stack_read_MUX[uxn_opcodes_h_l1414_c7_1a71] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;

     -- t8_MUX[uxn_opcodes_h_l1414_c7_1a71] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1414_c7_1a71_cond <= VAR_t8_MUX_uxn_opcodes_h_l1414_c7_1a71_cond;
     t8_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue;
     t8_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output := t8_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1426_c7_fc7f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1426_c7_fc7f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1420_c7_7f85] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1420_c7_7f85] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1418_c32_c41c] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_left;
     BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_return_output := BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1405_c1_246e] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1420_c7_7f85] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output := result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1418_c32_79e3_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1418_c32_c41c_return_output;
     VAR_printf_uxn_opcodes_h_l1406_c3_7745_uxn_opcodes_h_l1406_c3_7745_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1405_c1_246e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_fc7f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;
     -- t8_MUX[uxn_opcodes_h_l1411_c7_a63d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1411_c7_a63d_cond <= VAR_t8_MUX_uxn_opcodes_h_l1411_c7_a63d_cond;
     t8_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue;
     t8_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output := t8_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1414_c7_1a71] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output := result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1420_c7_7f85] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1414_c7_1a71] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1411_c7_a63d] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;

     -- printf_uxn_opcodes_h_l1406_c3_7745[uxn_opcodes_h_l1406_c3_7745] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1406_c3_7745_uxn_opcodes_h_l1406_c3_7745_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1406_c3_7745_uxn_opcodes_h_l1406_c3_7745_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1420_c7_7f85] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1414_c7_1a71] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;

     -- MUX[uxn_opcodes_h_l1418_c32_79e3] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1418_c32_79e3_cond <= VAR_MUX_uxn_opcodes_h_l1418_c32_79e3_cond;
     MUX_uxn_opcodes_h_l1418_c32_79e3_iftrue <= VAR_MUX_uxn_opcodes_h_l1418_c32_79e3_iftrue;
     MUX_uxn_opcodes_h_l1418_c32_79e3_iffalse <= VAR_MUX_uxn_opcodes_h_l1418_c32_79e3_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1418_c32_79e3_return_output := MUX_uxn_opcodes_h_l1418_c32_79e3_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue := VAR_MUX_uxn_opcodes_h_l1418_c32_79e3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1420_c7_7f85_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;
     -- result_is_stack_read_MUX[uxn_opcodes_h_l1405_c2_24aa] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1414_c7_1a71] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1414_c7_1a71] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;

     -- t8_MUX[uxn_opcodes_h_l1405_c2_24aa] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1405_c2_24aa_cond <= VAR_t8_MUX_uxn_opcodes_h_l1405_c2_24aa_cond;
     t8_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue;
     t8_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output := t8_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1411_c7_a63d] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output := result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1411_c7_a63d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1414_c7_1a71] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1411_c7_a63d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1414_c7_1a71_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1405_c2_24aa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1405_c2_24aa] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output := result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1411_c7_a63d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1405_c2_24aa] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1411_c7_a63d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1411_c7_a63d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1411_c7_a63d_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1405_c2_24aa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1405_c2_24aa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1405_c2_24aa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_28d7_uxn_opcodes_h_l1401_l1431_DUPLICATE_3816 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_28d7_uxn_opcodes_h_l1401_l1431_DUPLICATE_3816_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_28d7(
     result,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1405_c2_24aa_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_28d7_uxn_opcodes_h_l1401_l1431_DUPLICATE_3816_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_28d7_uxn_opcodes_h_l1401_l1431_DUPLICATE_3816_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
