-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity div_0CLK_4e24eea7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end div_0CLK_4e24eea7;
architecture arch of div_0CLK_4e24eea7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2056_c6_41f6]
signal BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2056_c2_135e]
signal result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2056_c2_135e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2056_c2_135e]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2056_c2_135e]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2056_c2_135e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2056_c2_135e]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2056_c2_135e]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2056_c2_135e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2056_c2_135e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2056_c2_135e]
signal t8_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2056_c2_135e]
signal n8_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2069_c11_b2cd]
signal BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2069_c7_5ef2]
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2069_c7_5ef2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2069_c7_5ef2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2069_c7_5ef2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2069_c7_5ef2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2069_c7_5ef2]
signal t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2069_c7_5ef2]
signal n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2072_c11_1025]
signal BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2072_c7_08af]
signal result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2072_c7_08af]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2072_c7_08af]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2072_c7_08af]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2072_c7_08af]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2072_c7_08af]
signal t8_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2072_c7_08af]
signal n8_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2075_c11_cb7f]
signal BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2075_c7_a7a9]
signal result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2075_c7_a7a9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2075_c7_a7a9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2075_c7_a7a9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2075_c7_a7a9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2075_c7_a7a9]
signal n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2077_c30_a6ff]
signal sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2080_c21_221f]
signal BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_return_output : unsigned(0 downto 0);

-- BIN_OP_DIV[uxn_opcodes_h_l2080_c35_469d]
signal BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_left : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_right : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l2080_c21_486f]
signal MUX_uxn_opcodes_h_l2080_c21_486f_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2080_c21_486f_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2080_c21_486f_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2080_c21_486f_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_243c( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : signed;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_pc_updated := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.sp_relative_shift := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6
BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_left,
BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_right,
BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_return_output);

-- t8_MUX_uxn_opcodes_h_l2056_c2_135e
t8_MUX_uxn_opcodes_h_l2056_c2_135e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2056_c2_135e_cond,
t8_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue,
t8_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse,
t8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output);

-- n8_MUX_uxn_opcodes_h_l2056_c2_135e
n8_MUX_uxn_opcodes_h_l2056_c2_135e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2056_c2_135e_cond,
n8_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue,
n8_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse,
n8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_left,
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_right,
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output);

-- t8_MUX_uxn_opcodes_h_l2069_c7_5ef2
t8_MUX_uxn_opcodes_h_l2069_c7_5ef2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond,
t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue,
t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse,
t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output);

-- n8_MUX_uxn_opcodes_h_l2069_c7_5ef2
n8_MUX_uxn_opcodes_h_l2069_c7_5ef2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond,
n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue,
n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse,
n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025
BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_left,
BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_right,
BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_cond,
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_return_output);

-- t8_MUX_uxn_opcodes_h_l2072_c7_08af
t8_MUX_uxn_opcodes_h_l2072_c7_08af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2072_c7_08af_cond,
t8_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue,
t8_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse,
t8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output);

-- n8_MUX_uxn_opcodes_h_l2072_c7_08af
n8_MUX_uxn_opcodes_h_l2072_c7_08af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2072_c7_08af_cond,
n8_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue,
n8_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse,
n8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f
BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_left,
BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_right,
BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond,
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output);

-- n8_MUX_uxn_opcodes_h_l2075_c7_a7a9
n8_MUX_uxn_opcodes_h_l2075_c7_a7a9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond,
n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue,
n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse,
n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff
sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_ins,
sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_x,
sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_y,
sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f
BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_left,
BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_right,
BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_return_output);

-- BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d
BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d : entity work.BIN_OP_DIV_uint8_t_uint8_t_0CLK_371b3c10 port map (
BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_left,
BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_right,
BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_return_output);

-- MUX_uxn_opcodes_h_l2080_c21_486f
MUX_uxn_opcodes_h_l2080_c21_486f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2080_c21_486f_cond,
MUX_uxn_opcodes_h_l2080_c21_486f_iftrue,
MUX_uxn_opcodes_h_l2080_c21_486f_iffalse,
MUX_uxn_opcodes_h_l2080_c21_486f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
 t8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
 n8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output,
 t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output,
 n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_return_output,
 t8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output,
 n8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output,
 n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output,
 sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_return_output,
 BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_return_output,
 MUX_uxn_opcodes_h_l2080_c21_486f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2066_c3_787c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2061_c3_46a5 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2056_c2_135e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2070_c3_bedf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2072_c7_08af_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2079_c3_1c5f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2080_c21_486f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2080_c21_486f_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2080_c21_486f_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2080_c21_486f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2072_l2056_l2075_l2069_DUPLICATE_ea75_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_b079_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_db81_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_614e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_89a3_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2084_l2052_DUPLICATE_16ec_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2079_c3_1c5f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2079_c3_1c5f;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2066_c3_787c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2066_c3_787c;
     VAR_MUX_uxn_opcodes_h_l2080_c21_486f_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2070_c3_bedf := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2070_c3_bedf;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_right := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2061_c3_46a5 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2061_c3_46a5;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_left := VAR_phase;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_right := t8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2075_c11_cb7f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2080_c21_221f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_614e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_614e_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2069_c11_b2cd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2077_c30_a6ff] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_ins;
     sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_x;
     sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_return_output := sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2056_c2_135e_return_output := result.is_vram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_db81 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_db81_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_89a3 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_89a3_return_output := result.stack_address_sp_offset;

     -- BIN_OP_DIV[uxn_opcodes_h_l2080_c35_469d] LATENCY=0
     -- Inputs
     BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_left <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_left;
     BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_right <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_right;
     -- Outputs
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_return_output := BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2072_l2056_l2075_l2069_DUPLICATE_ea75 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2072_l2056_l2075_l2069_DUPLICATE_ea75_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2072_c11_1025] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_left;
     BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_return_output := BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2056_c2_135e_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2056_c6_41f6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2056_c2_135e_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_b079 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_b079_return_output := result.is_stack_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2056_c2_135e_return_output := result.is_pc_updated;

     -- Submodule level 1
     VAR_MUX_uxn_opcodes_h_l2080_c21_486f_iffalse := VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_469d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2056_c2_135e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2056_c2_135e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_41f6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_b2cd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2072_c7_08af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2072_c7_08af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_1025_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_cb7f_return_output;
     VAR_MUX_uxn_opcodes_h_l2080_c21_486f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_221f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_db81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_db81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_db81_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_614e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_614e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_614e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_b079_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_b079_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2072_l2075_l2069_DUPLICATE_b079_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_89a3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_89a3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2072_l2056_l2075_l2069_DUPLICATE_ea75_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2072_l2056_l2075_l2069_DUPLICATE_ea75_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2072_l2056_l2075_l2069_DUPLICATE_ea75_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2072_l2056_l2075_l2069_DUPLICATE_ea75_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2056_c2_135e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2056_c2_135e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2056_c2_135e_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2056_c2_135e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_a6ff_return_output;
     -- t8_MUX[uxn_opcodes_h_l2072_c7_08af] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2072_c7_08af_cond <= VAR_t8_MUX_uxn_opcodes_h_l2072_c7_08af_cond;
     t8_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue;
     t8_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output := t8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2075_c7_a7a9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output;

     -- MUX[uxn_opcodes_h_l2080_c21_486f] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2080_c21_486f_cond <= VAR_MUX_uxn_opcodes_h_l2080_c21_486f_cond;
     MUX_uxn_opcodes_h_l2080_c21_486f_iftrue <= VAR_MUX_uxn_opcodes_h_l2080_c21_486f_iftrue;
     MUX_uxn_opcodes_h_l2080_c21_486f_iffalse <= VAR_MUX_uxn_opcodes_h_l2080_c21_486f_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2080_c21_486f_return_output := MUX_uxn_opcodes_h_l2080_c21_486f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2075_c7_a7a9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output;

     -- n8_MUX[uxn_opcodes_h_l2075_c7_a7a9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond <= VAR_n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond;
     n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue;
     n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output := n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2075_c7_a7a9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2075_c7_a7a9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue := VAR_MUX_uxn_opcodes_h_l2080_c21_486f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;
     -- n8_MUX[uxn_opcodes_h_l2072_c7_08af] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2072_c7_08af_cond <= VAR_n8_MUX_uxn_opcodes_h_l2072_c7_08af_cond;
     n8_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue;
     n8_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output := n8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2072_c7_08af] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;

     -- t8_MUX[uxn_opcodes_h_l2069_c7_5ef2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond <= VAR_t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond;
     t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue;
     t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output := t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2072_c7_08af] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2072_c7_08af] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2075_c7_a7a9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output := result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2072_c7_08af] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_a7a9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2069_c7_5ef2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;

     -- t8_MUX[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2056_c2_135e_cond <= VAR_t8_MUX_uxn_opcodes_h_l2056_c2_135e_cond;
     t8_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue;
     t8_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output := t8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2072_c7_08af] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_return_output := result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2069_c7_5ef2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2069_c7_5ef2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;

     -- n8_MUX[uxn_opcodes_h_l2069_c7_5ef2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond <= VAR_n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond;
     n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue;
     n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output := n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2069_c7_5ef2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_08af_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2069_c7_5ef2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2056_c2_135e_cond <= VAR_n8_MUX_uxn_opcodes_h_l2056_c2_135e_cond;
     n8_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue;
     n8_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output := n8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2056_c2_135e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_5ef2_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2056_c2_135e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2084_l2052_DUPLICATE_16ec LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2084_l2052_DUPLICATE_16ec_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_243c(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_135e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_135e_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2084_l2052_DUPLICATE_16ec_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2084_l2052_DUPLICATE_16ec_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
