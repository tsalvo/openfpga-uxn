-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 43
entity inc_0CLK_66ba3dc0 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc_0CLK_66ba3dc0;
architecture arch of inc_0CLK_66ba3dc0 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1527_c6_7e5d]
signal BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1527_c1_f775]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1527_c2_c788]
signal t8_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1527_c2_c788]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1527_c2_c788]
signal result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1527_c2_c788]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1527_c2_c788]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : signed(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1527_c2_c788]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1527_c2_c788]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1527_c2_c788]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l1528_c3_ea7f[uxn_opcodes_h_l1528_c3_ea7f]
signal printf_uxn_opcodes_h_l1528_c3_ea7f_uxn_opcodes_h_l1528_c3_ea7f_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1533_c11_71b1]
signal BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1533_c7_f956]
signal t8_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1533_c7_f956]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1533_c7_f956]
signal result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1533_c7_f956]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1533_c7_f956]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : signed(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1533_c7_f956]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1533_c7_f956]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1533_c7_f956]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1536_c11_6e3c]
signal BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1536_c7_efeb]
signal t8_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1536_c7_efeb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1536_c7_efeb]
signal result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1536_c7_efeb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1536_c7_efeb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : signed(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1536_c7_efeb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1536_c7_efeb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1536_c7_efeb]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1540_c32_8469]
signal BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1540_c32_4919]
signal BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1540_c32_d13e]
signal MUX_uxn_opcodes_h_l1540_c32_d13e_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1540_c32_d13e_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1540_c32_d13e_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1540_c32_d13e_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1542_c11_ca7a]
signal BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1542_c7_7c6b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1542_c7_7c6b]
signal result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1542_c7_7c6b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1542_c7_7c6b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1542_c7_7c6b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1546_c24_6eb0]
signal BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1548_c11_080d]
signal BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1548_c7_c2e5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1548_c7_c2e5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_287e( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_sp_shift := ref_toks_1;
      base.stack_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.is_stack_read := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d
BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_left,
BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_right,
BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_return_output);

-- t8_MUX_uxn_opcodes_h_l1527_c2_c788
t8_MUX_uxn_opcodes_h_l1527_c2_c788 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1527_c2_c788_cond,
t8_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue,
t8_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse,
t8_MUX_uxn_opcodes_h_l1527_c2_c788_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788
result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788
result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_cond,
result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788
result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788
result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788
result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788
result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_return_output);

-- printf_uxn_opcodes_h_l1528_c3_ea7f_uxn_opcodes_h_l1528_c3_ea7f
printf_uxn_opcodes_h_l1528_c3_ea7f_uxn_opcodes_h_l1528_c3_ea7f : entity work.printf_uxn_opcodes_h_l1528_c3_ea7f_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1528_c3_ea7f_uxn_opcodes_h_l1528_c3_ea7f_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1
BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_left,
BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_right,
BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output);

-- t8_MUX_uxn_opcodes_h_l1533_c7_f956
t8_MUX_uxn_opcodes_h_l1533_c7_f956 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1533_c7_f956_cond,
t8_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue,
t8_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse,
t8_MUX_uxn_opcodes_h_l1533_c7_f956_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956
result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956
result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_cond,
result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956
result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956
result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956
result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956
result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c
BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_left,
BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_right,
BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output);

-- t8_MUX_uxn_opcodes_h_l1536_c7_efeb
t8_MUX_uxn_opcodes_h_l1536_c7_efeb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1536_c7_efeb_cond,
t8_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue,
t8_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse,
t8_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb
result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb
result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_cond,
result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb
result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb
result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb
result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb
result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469
BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_left,
BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_right,
BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919
BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_left,
BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_right,
BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_return_output);

-- MUX_uxn_opcodes_h_l1540_c32_d13e
MUX_uxn_opcodes_h_l1540_c32_d13e : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1540_c32_d13e_cond,
MUX_uxn_opcodes_h_l1540_c32_d13e_iftrue,
MUX_uxn_opcodes_h_l1540_c32_d13e_iffalse,
MUX_uxn_opcodes_h_l1540_c32_d13e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a
BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_left,
BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_right,
BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b
result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b
result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond,
result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b
result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b
result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0
BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_left,
BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_right,
BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d
BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_left,
BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_right,
BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5
result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5
result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_return_output,
 t8_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output,
 t8_MUX_uxn_opcodes_h_l1533_c7_f956_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output,
 t8_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_return_output,
 MUX_uxn_opcodes_h_l1540_c32_d13e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1530_c3_8d79 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1528_c3_ea7f_uxn_opcodes_h_l1528_c3_ea7f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1534_c3_053e : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1540_c32_d13e_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1540_c32_d13e_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1540_c32_d13e_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1540_c32_d13e_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_uxn_opcodes_h_l1546_c3_ed88 : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1545_c3_63d4 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_return_output : unsigned(8 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1527_l1542_l1533_DUPLICATE_f807_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1527_l1542_l1533_l1536_DUPLICATE_650e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1527_l1533_l1548_l1536_DUPLICATE_9c89_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1527_l1533_l1536_DUPLICATE_61a3_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1542_l1533_l1548_l1536_DUPLICATE_5852_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1533_l1536_DUPLICATE_bac0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1542_l1536_DUPLICATE_38f3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_287e_uxn_opcodes_h_l1553_l1523_DUPLICATE_b237_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_right := to_unsigned(0, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_right := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_right := to_unsigned(128, 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1534_c3_053e := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1534_c3_053e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1545_c3_63d4 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1545_c3_63d4;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1540_c32_d13e_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_MUX_uxn_opcodes_h_l1540_c32_d13e_iffalse := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1530_c3_8d79 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1530_c3_8d79;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1542_l1533_l1548_l1536_DUPLICATE_5852 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1542_l1533_l1548_l1536_DUPLICATE_5852_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1548_c11_080d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1527_c6_7e5d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1533_l1536_DUPLICATE_bac0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1533_l1536_DUPLICATE_bac0_return_output := result.is_stack_read;

     -- BIN_OP_EQ[uxn_opcodes_h_l1542_c11_ca7a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1536_c11_6e3c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1546_c24_6eb0] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1527_l1542_l1533_DUPLICATE_f807 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1527_l1542_l1533_DUPLICATE_f807_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1533_c11_71b1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l1540_c32_8469] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_left;
     BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_return_output := BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1542_l1536_DUPLICATE_38f3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1542_l1536_DUPLICATE_38f3_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1527_l1533_l1536_DUPLICATE_61a3 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1527_l1533_l1536_DUPLICATE_61a3_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1527_l1542_l1533_l1536_DUPLICATE_650e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1527_l1542_l1533_l1536_DUPLICATE_650e_return_output := result.stack_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1527_l1533_l1548_l1536_DUPLICATE_9c89 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1527_l1533_l1548_l1536_DUPLICATE_9c89_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1540_c32_8469_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1527_c2_c788_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1527_c6_7e5d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1533_c7_f956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1533_c11_71b1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1536_c7_efeb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_6e3c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_ca7a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1548_c11_080d_return_output;
     VAR_result_stack_value_uxn_opcodes_h_l1546_c3_ed88 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1546_c24_6eb0_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1527_l1533_l1536_DUPLICATE_61a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1527_l1533_l1536_DUPLICATE_61a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1527_l1533_l1536_DUPLICATE_61a3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1542_l1533_l1548_l1536_DUPLICATE_5852_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1542_l1533_l1548_l1536_DUPLICATE_5852_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1542_l1533_l1548_l1536_DUPLICATE_5852_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1542_l1533_l1548_l1536_DUPLICATE_5852_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1527_l1542_l1533_DUPLICATE_f807_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1527_l1542_l1533_DUPLICATE_f807_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1527_l1542_l1533_DUPLICATE_f807_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1533_l1536_DUPLICATE_bac0_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1533_l1536_DUPLICATE_bac0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1527_l1533_l1548_l1536_DUPLICATE_9c89_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1527_l1533_l1548_l1536_DUPLICATE_9c89_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1527_l1533_l1548_l1536_DUPLICATE_9c89_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1527_l1533_l1548_l1536_DUPLICATE_9c89_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1542_l1536_DUPLICATE_38f3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1542_l1536_DUPLICATE_38f3_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1527_l1542_l1533_l1536_DUPLICATE_650e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1527_l1542_l1533_l1536_DUPLICATE_650e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1527_l1542_l1533_l1536_DUPLICATE_650e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1527_l1542_l1533_l1536_DUPLICATE_650e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue := VAR_result_stack_value_uxn_opcodes_h_l1546_c3_ed88;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1542_c7_7c6b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1536_c7_efeb] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1536_c7_efeb_cond <= VAR_t8_MUX_uxn_opcodes_h_l1536_c7_efeb_cond;
     t8_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue;
     t8_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output := t8_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1542_c7_7c6b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1536_c7_efeb] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1527_c1_f775] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1540_c32_4919] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_left;
     BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_return_output := BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1542_c7_7c6b] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output := result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1548_c7_c2e5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1548_c7_c2e5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1540_c32_d13e_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1540_c32_4919_return_output;
     VAR_printf_uxn_opcodes_h_l1528_c3_ea7f_uxn_opcodes_h_l1528_c3_ea7f_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1527_c1_f775_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1548_c7_c2e5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1542_c7_7c6b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output;

     -- printf_uxn_opcodes_h_l1528_c3_ea7f[uxn_opcodes_h_l1528_c3_ea7f] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1528_c3_ea7f_uxn_opcodes_h_l1528_c3_ea7f_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1528_c3_ea7f_uxn_opcodes_h_l1528_c3_ea7f_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- t8_MUX[uxn_opcodes_h_l1533_c7_f956] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1533_c7_f956_cond <= VAR_t8_MUX_uxn_opcodes_h_l1533_c7_f956_cond;
     t8_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue;
     t8_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1533_c7_f956_return_output := t8_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1533_c7_f956] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1536_c7_efeb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1542_c7_7c6b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1536_c7_efeb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;

     -- MUX[uxn_opcodes_h_l1540_c32_d13e] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1540_c32_d13e_cond <= VAR_MUX_uxn_opcodes_h_l1540_c32_d13e_cond;
     MUX_uxn_opcodes_h_l1540_c32_d13e_iftrue <= VAR_MUX_uxn_opcodes_h_l1540_c32_d13e_iftrue;
     MUX_uxn_opcodes_h_l1540_c32_d13e_iffalse <= VAR_MUX_uxn_opcodes_h_l1540_c32_d13e_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1540_c32_d13e_return_output := MUX_uxn_opcodes_h_l1540_c32_d13e_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1536_c7_efeb] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output := result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue := VAR_MUX_uxn_opcodes_h_l1540_c32_d13e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_7c6b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;
     -- result_stack_value_MUX[uxn_opcodes_h_l1533_c7_f956] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_return_output := result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1527_c2_c788] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1536_c7_efeb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;

     -- t8_MUX[uxn_opcodes_h_l1527_c2_c788] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1527_c2_c788_cond <= VAR_t8_MUX_uxn_opcodes_h_l1527_c2_c788_cond;
     t8_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue;
     t8_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1527_c2_c788_return_output := t8_MUX_uxn_opcodes_h_l1527_c2_c788_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1536_c7_efeb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1533_c7_f956] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1536_c7_efeb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1533_c7_f956] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1536_c7_efeb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1527_c2_c788_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1533_c7_f956] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1533_c7_f956] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1527_c2_c788] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1527_c2_c788] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_return_output := result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1533_c7_f956] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1527_c2_c788] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1533_c7_f956_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1527_c2_c788] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1527_c2_c788] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1527_c2_c788] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_287e_uxn_opcodes_h_l1553_l1523_DUPLICATE_b237 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_287e_uxn_opcodes_h_l1553_l1523_DUPLICATE_b237_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_287e(
     result,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1527_c2_c788_return_output,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1527_c2_c788_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_287e_uxn_opcodes_h_l1553_l1523_DUPLICATE_b237_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_287e_uxn_opcodes_h_l1553_l1523_DUPLICATE_b237_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
