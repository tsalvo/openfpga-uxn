-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 43
entity inc_0CLK_66ba3dc0 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc_0CLK_66ba3dc0;
architecture arch of inc_0CLK_66ba3dc0 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(15 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1030_c6_8914]
signal BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1030_c1_770e]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1030_c2_fb7e]
signal t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(15 downto 0);
signal t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(15 downto 0);
signal t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(15 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1030_c2_fb7e]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1030_c2_fb7e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1030_c2_fb7e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1030_c2_fb7e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1030_c2_fb7e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1030_c2_fb7e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1030_c2_fb7e]
signal result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1031_c3_a87d[uxn_opcodes_h_l1031_c3_a87d]
signal printf_uxn_opcodes_h_l1031_c3_a87d_uxn_opcodes_h_l1031_c3_a87d_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1036_c11_d92b]
signal BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1036_c7_3a4f]
signal t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(15 downto 0);
signal t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(15 downto 0);
signal t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(15 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1036_c7_3a4f]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1036_c7_3a4f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1036_c7_3a4f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1036_c7_3a4f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1036_c7_3a4f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1036_c7_3a4f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1036_c7_3a4f]
signal result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1039_c11_6202]
signal BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1039_c7_0368]
signal t8_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(15 downto 0);
signal t8_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(15 downto 0);
signal t8_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(15 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l1039_c7_0368]
signal result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1039_c7_0368]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : signed(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1039_c7_0368]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1039_c7_0368]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1039_c7_0368]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1039_c7_0368]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1039_c7_0368]
signal result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(7 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1043_c32_57be]
signal BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1043_c32_9bf5]
signal BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1043_c32_5c83]
signal MUX_uxn_opcodes_h_l1043_c32_5c83_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1043_c32_5c83_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1043_c32_5c83_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1043_c32_5c83_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1045_c11_289a]
signal BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1045_c7_db6f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1045_c7_db6f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1045_c7_db6f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1045_c7_db6f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1045_c7_db6f]
signal result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1049_c24_9ad1]
signal BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1051_c11_976c]
signal BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1051_c7_f08a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1051_c7_f08a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_28d7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : signed;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_read := ref_toks_1;
      base.sp_relative_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_sp_shift := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.stack_value := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914
BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_left,
BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_right,
BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_return_output);

-- t8_MUX_uxn_opcodes_h_l1030_c2_fb7e
t8_MUX_uxn_opcodes_h_l1030_c2_fb7e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond,
t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue,
t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse,
t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e
result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e
result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e
result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e
result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e
result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond,
result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output);

-- printf_uxn_opcodes_h_l1031_c3_a87d_uxn_opcodes_h_l1031_c3_a87d
printf_uxn_opcodes_h_l1031_c3_a87d_uxn_opcodes_h_l1031_c3_a87d : entity work.printf_uxn_opcodes_h_l1031_c3_a87d_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1031_c3_a87d_uxn_opcodes_h_l1031_c3_a87d_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b
BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_left,
BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_right,
BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output);

-- t8_MUX_uxn_opcodes_h_l1036_c7_3a4f
t8_MUX_uxn_opcodes_h_l1036_c7_3a4f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond,
t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue,
t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse,
t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f
result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f
result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f
result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f
result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f
result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond,
result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202
BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_left,
BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_right,
BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output);

-- t8_MUX_uxn_opcodes_h_l1039_c7_0368
t8_MUX_uxn_opcodes_h_l1039_c7_0368 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1039_c7_0368_cond,
t8_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue,
t8_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse,
t8_MUX_uxn_opcodes_h_l1039_c7_0368_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368
result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368
result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368
result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368
result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368
result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368
result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_cond,
result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be
BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_left,
BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_right,
BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5
BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_left,
BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_right,
BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_return_output);

-- MUX_uxn_opcodes_h_l1043_c32_5c83
MUX_uxn_opcodes_h_l1043_c32_5c83 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1043_c32_5c83_cond,
MUX_uxn_opcodes_h_l1043_c32_5c83_iftrue,
MUX_uxn_opcodes_h_l1043_c32_5c83_iffalse,
MUX_uxn_opcodes_h_l1043_c32_5c83_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a
BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_left,
BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_right,
BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f
result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f
result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f
result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f
result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_cond,
result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1
BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1 : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_left,
BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_right,
BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c
BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_left,
BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_right,
BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a
result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a
result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_return_output,
 t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output,
 t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output,
 t8_MUX_uxn_opcodes_h_l1039_c7_0368_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_return_output,
 MUX_uxn_opcodes_h_l1043_c32_5c83_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1033_c3_9700 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1031_c3_a87d_uxn_opcodes_h_l1031_c3_a87d_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1037_c3_dfa9 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(15 downto 0);
 variable VAR_t8_uxn_opcodes_h_l1040_c3_366c : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(15 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1043_c32_5c83_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1043_c32_5c83_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1043_c32_5c83_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1043_c32_5c83_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1048_c3_a93f : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_uxn_opcodes_h_l1049_c3_ced6 : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1036_l1039_l1030_DUPLICATE_8d1c_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1030_DUPLICATE_1c66_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1036_l1030_l1045_DUPLICATE_c30c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1036_l1039_l1030_l1045_DUPLICATE_561c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1036_l1039_DUPLICATE_6bc5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1045_DUPLICATE_a56d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1039_l1045_DUPLICATE_d533_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_28d7_uxn_opcodes_h_l1026_l1056_DUPLICATE_54fd_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(15 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1048_c3_a93f := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1048_c3_a93f;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1043_c32_5c83_iffalse := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_right := to_unsigned(2, 2);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1043_c32_5c83_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1037_c3_dfa9 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1037_c3_dfa9;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_right := to_unsigned(1, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_right := to_unsigned(128, 8);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1033_c3_9700 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1033_c3_9700;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_right := to_unsigned(4, 3);
     VAR_BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_left := VAR_phase;
     VAR_t8_uxn_opcodes_h_l1040_c3_366c := resize(VAR_previous_stack_read, 16);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse := t8;
     REG_VAR_tmp16 := tmp16;
     VAR_t8_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue := VAR_t8_uxn_opcodes_h_l1040_c3_366c;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1036_l1039_DUPLICATE_6bc5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1036_l1039_DUPLICATE_6bc5_return_output := result.is_stack_read;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1036_l1030_l1045_DUPLICATE_c30c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1036_l1030_l1045_DUPLICATE_c30c_return_output := result.is_sp_shift;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1036_l1039_l1030_DUPLICATE_8d1c LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1036_l1039_l1030_DUPLICATE_8d1c_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1039_l1045_DUPLICATE_d533 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1039_l1045_DUPLICATE_d533_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1045_DUPLICATE_a56d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1045_DUPLICATE_a56d_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1036_l1039_l1030_l1045_DUPLICATE_561c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1036_l1039_l1030_l1045_DUPLICATE_561c_return_output := result.stack_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1030_DUPLICATE_1c66 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1030_DUPLICATE_1c66_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1045_c11_289a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1036_c11_d92b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1039_c11_6202] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_left;
     BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output := BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1030_c6_8914] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_left;
     BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output := BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1049_c24_9ad1] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1051_c11_976c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l1043_c32_57be] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_left;
     BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_return_output := BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1043_c32_57be_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1030_c6_8914_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1036_c11_d92b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1039_c7_0368_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_6202_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c11_289a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_976c_return_output;
     VAR_result_stack_value_uxn_opcodes_h_l1049_c3_ced6 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1049_c24_9ad1_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1036_l1039_l1030_DUPLICATE_8d1c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1036_l1039_l1030_DUPLICATE_8d1c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1036_l1039_l1030_DUPLICATE_8d1c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1045_DUPLICATE_a56d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1045_DUPLICATE_a56d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1045_DUPLICATE_a56d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1045_DUPLICATE_a56d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1036_l1030_l1045_DUPLICATE_c30c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1036_l1030_l1045_DUPLICATE_c30c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1036_l1030_l1045_DUPLICATE_c30c_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1036_l1039_DUPLICATE_6bc5_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l1036_l1039_DUPLICATE_6bc5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1030_DUPLICATE_1c66_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1030_DUPLICATE_1c66_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1030_DUPLICATE_1c66_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1036_l1051_l1039_l1030_DUPLICATE_1c66_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1039_l1045_DUPLICATE_d533_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1039_l1045_DUPLICATE_d533_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1036_l1039_l1030_l1045_DUPLICATE_561c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1036_l1039_l1030_l1045_DUPLICATE_561c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1036_l1039_l1030_l1045_DUPLICATE_561c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1036_l1039_l1030_l1045_DUPLICATE_561c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue := VAR_result_stack_value_uxn_opcodes_h_l1049_c3_ced6;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1051_c7_f08a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1051_c7_f08a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1043_c32_9bf5] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_left;
     BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_return_output := BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1039_c7_0368] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;

     -- t8_MUX[uxn_opcodes_h_l1039_c7_0368] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1039_c7_0368_cond <= VAR_t8_MUX_uxn_opcodes_h_l1039_c7_0368_cond;
     t8_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue;
     t8_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1039_c7_0368_return_output := t8_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1030_c1_770e] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1045_c7_db6f] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output := result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1045_c7_db6f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1045_c7_db6f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1043_c32_5c83_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1043_c32_9bf5_return_output;
     VAR_printf_uxn_opcodes_h_l1031_c3_a87d_uxn_opcodes_h_l1031_c3_a87d_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1030_c1_770e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_f08a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;
     -- result_is_stack_read_MUX[uxn_opcodes_h_l1036_c7_3a4f] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1045_c7_db6f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1039_c7_0368] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_return_output := result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1039_c7_0368] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;

     -- MUX[uxn_opcodes_h_l1043_c32_5c83] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1043_c32_5c83_cond <= VAR_MUX_uxn_opcodes_h_l1043_c32_5c83_cond;
     MUX_uxn_opcodes_h_l1043_c32_5c83_iftrue <= VAR_MUX_uxn_opcodes_h_l1043_c32_5c83_iftrue;
     MUX_uxn_opcodes_h_l1043_c32_5c83_iffalse <= VAR_MUX_uxn_opcodes_h_l1043_c32_5c83_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1043_c32_5c83_return_output := MUX_uxn_opcodes_h_l1043_c32_5c83_return_output;

     -- printf_uxn_opcodes_h_l1031_c3_a87d[uxn_opcodes_h_l1031_c3_a87d] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1031_c3_a87d_uxn_opcodes_h_l1031_c3_a87d_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1031_c3_a87d_uxn_opcodes_h_l1031_c3_a87d_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1039_c7_0368] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1045_c7_db6f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1036_c7_3a4f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond;
     t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue;
     t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output := t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue := VAR_MUX_uxn_opcodes_h_l1043_c32_5c83_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c7_db6f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;
     -- t8_MUX[uxn_opcodes_h_l1030_c2_fb7e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond <= VAR_t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond;
     t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue;
     t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output := t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1036_c7_3a4f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1039_c7_0368] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1036_c7_3a4f] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output := result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1036_c7_3a4f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l1030_c2_fb7e] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1039_c7_0368] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1039_c7_0368] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1039_c7_0368_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1036_c7_3a4f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1036_c7_3a4f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1036_c7_3a4f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1030_c2_fb7e] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output := result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1030_c2_fb7e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1030_c2_fb7e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1036_c7_3a4f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1030_c2_fb7e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1030_c2_fb7e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1030_c2_fb7e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_28d7_uxn_opcodes_h_l1026_l1056_DUPLICATE_54fd LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_28d7_uxn_opcodes_h_l1026_l1056_DUPLICATE_54fd_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_28d7(
     result,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1030_c2_fb7e_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_28d7_uxn_opcodes_h_l1026_l1056_DUPLICATE_54fd_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_28d7_uxn_opcodes_h_l1026_l1056_DUPLICATE_54fd_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
