-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity jcn_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jcn_0CLK_f62d646e;
architecture arch of jcn_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l688_c6_4aef]
signal BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l688_c2_e9c3]
signal n8_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l688_c2_e9c3]
signal t8_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l688_c2_e9c3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l688_c2_e9c3]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l688_c2_e9c3]
signal result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l688_c2_e9c3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l688_c2_e9c3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l688_c2_e9c3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l693_c11_ee9f]
signal BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l693_c7_d654]
signal n8_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l693_c7_d654]
signal t8_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l693_c7_d654]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l693_c7_d654]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l693_c7_d654]
signal result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l693_c7_d654]
signal result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l693_c7_d654]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l693_c7_d654]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l696_c11_2f95]
signal BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l696_c7_1244]
signal n8_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l696_c7_1244]
signal t8_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l696_c7_1244]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l696_c7_1244]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l696_c7_1244]
signal result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l696_c7_1244]
signal result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l696_c7_1244]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l696_c7_1244]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l700_c11_902c]
signal BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l700_c7_c6fe]
signal n8_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l700_c7_c6fe]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l700_c7_c6fe]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l700_c7_c6fe]
signal result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l700_c7_c6fe]
signal result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l700_c7_c6fe]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l700_c7_c6fe]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l703_c11_d614]
signal BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l703_c7_a5f9]
signal n8_MUX_uxn_opcodes_h_l703_c7_a5f9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l703_c7_a5f9]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l703_c7_a5f9]
signal result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l703_c7_a5f9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l703_c7_a5f9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l703_c7_a5f9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l706_c30_e380]
signal sp_relative_shift_uxn_opcodes_h_l706_c30_e380_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l706_c30_e380_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l706_c30_e380_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l706_c30_e380_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l708_c22_4b6d]
signal BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l708_c37_c0c6]
signal BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_return_output : signed(17 downto 0);

-- MUX[uxn_opcodes_h_l708_c22_25d4]
signal MUX_uxn_opcodes_h_l708_c22_25d4_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l708_c22_25d4_iftrue : unsigned(15 downto 0);
signal MUX_uxn_opcodes_h_l708_c22_25d4_iffalse : unsigned(15 downto 0);
signal MUX_uxn_opcodes_h_l708_c22_25d4_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l710_c11_d691]
signal BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l710_c7_cb4c]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l710_c7_cb4c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l710_c7_cb4c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef
BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_left,
BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_right,
BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output);

-- n8_MUX_uxn_opcodes_h_l688_c2_e9c3
n8_MUX_uxn_opcodes_h_l688_c2_e9c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l688_c2_e9c3_cond,
n8_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue,
n8_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse,
n8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output);

-- t8_MUX_uxn_opcodes_h_l688_c2_e9c3
t8_MUX_uxn_opcodes_h_l688_c2_e9c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l688_c2_e9c3_cond,
t8_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue,
t8_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse,
t8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3
result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3
result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_cond,
result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3
result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3
result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3
result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f
BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_left,
BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_right,
BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output);

-- n8_MUX_uxn_opcodes_h_l693_c7_d654
n8_MUX_uxn_opcodes_h_l693_c7_d654 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l693_c7_d654_cond,
n8_MUX_uxn_opcodes_h_l693_c7_d654_iftrue,
n8_MUX_uxn_opcodes_h_l693_c7_d654_iffalse,
n8_MUX_uxn_opcodes_h_l693_c7_d654_return_output);

-- t8_MUX_uxn_opcodes_h_l693_c7_d654
t8_MUX_uxn_opcodes_h_l693_c7_d654 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l693_c7_d654_cond,
t8_MUX_uxn_opcodes_h_l693_c7_d654_iftrue,
t8_MUX_uxn_opcodes_h_l693_c7_d654_iffalse,
t8_MUX_uxn_opcodes_h_l693_c7_d654_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654
result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654
result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_cond,
result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654
result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654
result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654
result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95
BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_left,
BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_right,
BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output);

-- n8_MUX_uxn_opcodes_h_l696_c7_1244
n8_MUX_uxn_opcodes_h_l696_c7_1244 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l696_c7_1244_cond,
n8_MUX_uxn_opcodes_h_l696_c7_1244_iftrue,
n8_MUX_uxn_opcodes_h_l696_c7_1244_iffalse,
n8_MUX_uxn_opcodes_h_l696_c7_1244_return_output);

-- t8_MUX_uxn_opcodes_h_l696_c7_1244
t8_MUX_uxn_opcodes_h_l696_c7_1244 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l696_c7_1244_cond,
t8_MUX_uxn_opcodes_h_l696_c7_1244_iftrue,
t8_MUX_uxn_opcodes_h_l696_c7_1244_iffalse,
t8_MUX_uxn_opcodes_h_l696_c7_1244_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244
result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244
result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_cond,
result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244
result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244
result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244
result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c
BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_left,
BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_right,
BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_return_output);

-- n8_MUX_uxn_opcodes_h_l700_c7_c6fe
n8_MUX_uxn_opcodes_h_l700_c7_c6fe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l700_c7_c6fe_cond,
n8_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue,
n8_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse,
n8_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe
result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe
result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_cond,
result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe
result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe
result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe
result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614
BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_left,
BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_right,
BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_return_output);

-- n8_MUX_uxn_opcodes_h_l703_c7_a5f9
n8_MUX_uxn_opcodes_h_l703_c7_a5f9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l703_c7_a5f9_cond,
n8_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue,
n8_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse,
n8_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9
result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9
result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_cond,
result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9
result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9
result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9
result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output);

-- sp_relative_shift_uxn_opcodes_h_l706_c30_e380
sp_relative_shift_uxn_opcodes_h_l706_c30_e380 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l706_c30_e380_ins,
sp_relative_shift_uxn_opcodes_h_l706_c30_e380_x,
sp_relative_shift_uxn_opcodes_h_l706_c30_e380_y,
sp_relative_shift_uxn_opcodes_h_l706_c30_e380_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d
BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_left,
BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_right,
BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6
BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_left,
BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_right,
BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_return_output);

-- MUX_uxn_opcodes_h_l708_c22_25d4
MUX_uxn_opcodes_h_l708_c22_25d4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l708_c22_25d4_cond,
MUX_uxn_opcodes_h_l708_c22_25d4_iftrue,
MUX_uxn_opcodes_h_l708_c22_25d4_iffalse,
MUX_uxn_opcodes_h_l708_c22_25d4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691
BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_left,
BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_right,
BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c
result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c
result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c
result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output,
 n8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output,
 t8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output,
 n8_MUX_uxn_opcodes_h_l693_c7_d654_return_output,
 t8_MUX_uxn_opcodes_h_l693_c7_d654_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output,
 n8_MUX_uxn_opcodes_h_l696_c7_1244_return_output,
 t8_MUX_uxn_opcodes_h_l696_c7_1244_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_return_output,
 n8_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_return_output,
 n8_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output,
 sp_relative_shift_uxn_opcodes_h_l706_c30_e380_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_return_output,
 MUX_uxn_opcodes_h_l708_c22_25d4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l690_c3_c1eb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l694_c3_50fa : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l698_c3_5b52 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l701_c3_0d4f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l700_c7_c6fe_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l703_c7_a5f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l706_c30_e380_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l706_c30_e380_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l706_c30_e380_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l706_c30_e380_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l708_c22_25d4_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l708_c22_25d4_iftrue : unsigned(15 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l708_c22_25d4_iffalse : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l708_c42_f935_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_return_output : signed(17 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l708_c22_25d4_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_4b89_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_ff5e_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_4d81_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_5bc2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l693_l696_l710_l700_l703_DUPLICATE_dc2a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c_uxn_opcodes_h_l716_l684_DUPLICATE_0b5b_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l698_c3_5b52 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l698_c3_5b52;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l694_c3_50fa := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l694_c3_50fa;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l701_c3_0d4f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l701_c3_0d4f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l706_c30_e380_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l706_c30_e380_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l690_c3_c1eb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l690_c3_c1eb;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l706_c30_e380_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l693_c7_d654_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l696_c7_1244_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse := n8;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_MUX_uxn_opcodes_h_l708_c22_25d4_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l696_c7_1244_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l693_c7_d654_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l696_c7_1244_iffalse := t8;
     -- CAST_TO_int8_t[uxn_opcodes_h_l708_c42_f935] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l708_c42_f935_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_5bc2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_5bc2_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l703_c11_d614] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_left;
     BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_return_output := BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l693_l696_l710_l700_l703_DUPLICATE_dc2a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l693_l696_l710_l700_l703_DUPLICATE_dc2a_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_ff5e LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_ff5e_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l700_c11_902c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_left;
     BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_return_output := BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_4d81 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_4d81_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l708_c22_4b6d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_left;
     BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_return_output := BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l710_c11_d691] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_left;
     BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_return_output := BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l696_c11_2f95] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_left;
     BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output := BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l700_c7_c6fe] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l700_c7_c6fe_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l706_c30_e380] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l706_c30_e380_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l706_c30_e380_ins;
     sp_relative_shift_uxn_opcodes_h_l706_c30_e380_x <= VAR_sp_relative_shift_uxn_opcodes_h_l706_c30_e380_x;
     sp_relative_shift_uxn_opcodes_h_l706_c30_e380_y <= VAR_sp_relative_shift_uxn_opcodes_h_l706_c30_e380_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l706_c30_e380_return_output := sp_relative_shift_uxn_opcodes_h_l706_c30_e380_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_4b89 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_4b89_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l688_c6_4aef] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_left;
     BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output := BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l693_c11_ee9f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_left;
     BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output := BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l688_c2_e9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l688_c2_e9c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l688_c6_4aef_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l693_c7_d654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l693_c7_d654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l693_c11_ee9f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l696_c7_1244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l696_c7_1244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l696_c11_2f95_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l700_c7_c6fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c11_902c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l703_c7_a5f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l703_c11_d614_return_output;
     VAR_MUX_uxn_opcodes_h_l708_c22_25d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l708_c22_4b6d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l710_c11_d691_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l708_c42_f935_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_4d81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_4d81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_4d81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_4d81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_4d81_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_ff5e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_ff5e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_ff5e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_ff5e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l693_l696_l700_l688_l703_DUPLICATE_ff5e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l693_l696_l710_l700_l703_DUPLICATE_dc2a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l693_l696_l710_l700_l703_DUPLICATE_dc2a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l693_l696_l710_l700_l703_DUPLICATE_dc2a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l693_l696_l710_l700_l703_DUPLICATE_dc2a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l693_l696_l710_l700_l703_DUPLICATE_dc2a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_4b89_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_4b89_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_4b89_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_4b89_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_4b89_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_5bc2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_5bc2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_5bc2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_5bc2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l693_l696_l710_l700_l688_DUPLICATE_5bc2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l700_c7_c6fe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l706_c30_e380_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l700_c7_c6fe] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;

     -- t8_MUX[uxn_opcodes_h_l696_c7_1244] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l696_c7_1244_cond <= VAR_t8_MUX_uxn_opcodes_h_l696_c7_1244_cond;
     t8_MUX_uxn_opcodes_h_l696_c7_1244_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l696_c7_1244_iftrue;
     t8_MUX_uxn_opcodes_h_l696_c7_1244_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l696_c7_1244_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l696_c7_1244_return_output := t8_MUX_uxn_opcodes_h_l696_c7_1244_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l703_c7_a5f9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output;

     -- n8_MUX[uxn_opcodes_h_l703_c7_a5f9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l703_c7_a5f9_cond <= VAR_n8_MUX_uxn_opcodes_h_l703_c7_a5f9_cond;
     n8_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue;
     n8_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output := n8_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l710_c7_cb4c] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l710_c7_cb4c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l708_c37_c0c6] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_left;
     BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_return_output := BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l710_c7_cb4c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l708_c22_25d4_iffalse := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l708_c37_c0c6_return_output)),16);
     VAR_n8_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse := VAR_n8_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l710_c7_cb4c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l693_c7_d654_iffalse := VAR_t8_MUX_uxn_opcodes_h_l696_c7_1244_return_output;
     -- n8_MUX[uxn_opcodes_h_l700_c7_c6fe] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l700_c7_c6fe_cond <= VAR_n8_MUX_uxn_opcodes_h_l700_c7_c6fe_cond;
     n8_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue;
     n8_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output := n8_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l703_c7_a5f9] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output;

     -- MUX[uxn_opcodes_h_l708_c22_25d4] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l708_c22_25d4_cond <= VAR_MUX_uxn_opcodes_h_l708_c22_25d4_cond;
     MUX_uxn_opcodes_h_l708_c22_25d4_iftrue <= VAR_MUX_uxn_opcodes_h_l708_c22_25d4_iftrue;
     MUX_uxn_opcodes_h_l708_c22_25d4_iffalse <= VAR_MUX_uxn_opcodes_h_l708_c22_25d4_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l708_c22_25d4_return_output := MUX_uxn_opcodes_h_l708_c22_25d4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l700_c7_c6fe] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l703_c7_a5f9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l703_c7_a5f9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l696_c7_1244] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_return_output;

     -- t8_MUX[uxn_opcodes_h_l693_c7_d654] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l693_c7_d654_cond <= VAR_t8_MUX_uxn_opcodes_h_l693_c7_d654_cond;
     t8_MUX_uxn_opcodes_h_l693_c7_d654_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l693_c7_d654_iftrue;
     t8_MUX_uxn_opcodes_h_l693_c7_d654_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l693_c7_d654_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l693_c7_d654_return_output := t8_MUX_uxn_opcodes_h_l693_c7_d654_return_output;

     -- Submodule level 3
     VAR_result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue := VAR_MUX_uxn_opcodes_h_l708_c22_25d4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l696_c7_1244_iffalse := VAR_n8_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l696_c7_1244_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse := VAR_t8_MUX_uxn_opcodes_h_l693_c7_d654_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l703_c7_a5f9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output := result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l700_c7_c6fe] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l700_c7_c6fe] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l693_c7_d654] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l700_c7_c6fe] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;

     -- t8_MUX[uxn_opcodes_h_l688_c2_e9c3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l688_c2_e9c3_cond <= VAR_t8_MUX_uxn_opcodes_h_l688_c2_e9c3_cond;
     t8_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue;
     t8_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output := t8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l696_c7_1244] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output;

     -- n8_MUX[uxn_opcodes_h_l696_c7_1244] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l696_c7_1244_cond <= VAR_n8_MUX_uxn_opcodes_h_l696_c7_1244_cond;
     n8_MUX_uxn_opcodes_h_l696_c7_1244_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l696_c7_1244_iftrue;
     n8_MUX_uxn_opcodes_h_l696_c7_1244_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l696_c7_1244_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l696_c7_1244_return_output := n8_MUX_uxn_opcodes_h_l696_c7_1244_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l693_c7_d654_iffalse := VAR_n8_MUX_uxn_opcodes_h_l696_c7_1244_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l693_c7_d654_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l703_c7_a5f9_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l696_c7_1244] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l688_c2_e9c3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output;

     -- n8_MUX[uxn_opcodes_h_l693_c7_d654] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l693_c7_d654_cond <= VAR_n8_MUX_uxn_opcodes_h_l693_c7_d654_cond;
     n8_MUX_uxn_opcodes_h_l693_c7_d654_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l693_c7_d654_iftrue;
     n8_MUX_uxn_opcodes_h_l693_c7_d654_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l693_c7_d654_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l693_c7_d654_return_output := n8_MUX_uxn_opcodes_h_l693_c7_d654_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l700_c7_c6fe] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_cond;
     result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output := result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l696_c7_1244] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l693_c7_d654] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l696_c7_1244] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse := VAR_n8_MUX_uxn_opcodes_h_l693_c7_d654_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l696_c7_1244_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l696_c7_1244_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l696_c7_1244_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c7_c6fe_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l693_c7_d654] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l693_c7_d654] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l693_c7_d654] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l688_c2_e9c3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l696_c7_1244] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_cond;
     result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_return_output := result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_return_output;

     -- n8_MUX[uxn_opcodes_h_l688_c2_e9c3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l688_c2_e9c3_cond <= VAR_n8_MUX_uxn_opcodes_h_l688_c2_e9c3_cond;
     n8_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue;
     n8_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output := n8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l693_c7_d654_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l693_c7_d654_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l693_c7_d654_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l696_c7_1244_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l693_c7_d654] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_cond;
     result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_return_output := result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l688_c2_e9c3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l688_c2_e9c3] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l688_c2_e9c3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output;

     -- Submodule level 7
     VAR_result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l693_c7_d654_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l688_c2_e9c3] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_cond;
     result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output := result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c_uxn_opcodes_h_l716_l684_DUPLICATE_0b5b LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c_uxn_opcodes_h_l716_l684_DUPLICATE_0b5b_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l688_c2_e9c3_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c_uxn_opcodes_h_l716_l684_DUPLICATE_0b5b_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c_uxn_opcodes_h_l716_l684_DUPLICATE_0b5b_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
