-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity dup_0CLK_a148083c is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_a148083c;
architecture arch of dup_0CLK_a148083c is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2711_c6_84f5]
signal BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2711_c1_c79e]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2711_c2_e9a2]
signal t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2711_c2_e9a2]
signal result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2711_c2_e9a2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2711_c2_e9a2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2711_c2_e9a2]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2711_c2_e9a2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2711_c2_e9a2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2711_c2_e9a2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l2712_c3_9a46[uxn_opcodes_h_l2712_c3_9a46]
signal printf_uxn_opcodes_h_l2712_c3_9a46_uxn_opcodes_h_l2712_c3_9a46_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2717_c11_0f6c]
signal BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2717_c7_e289]
signal t8_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2717_c7_e289]
signal result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2717_c7_e289]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2717_c7_e289]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2717_c7_e289]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2717_c7_e289]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2717_c7_e289]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2717_c7_e289]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2720_c11_557b]
signal BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2720_c7_6f9b]
signal t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2720_c7_6f9b]
signal result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2720_c7_6f9b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2720_c7_6f9b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2720_c7_6f9b]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2720_c7_6f9b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2720_c7_6f9b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2720_c7_6f9b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2724_c32_ef56]
signal BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l2724_c32_c2a9]
signal BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l2724_c32_475a]
signal MUX_uxn_opcodes_h_l2724_c32_475a_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2724_c32_475a_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2724_c32_475a_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2724_c32_475a_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2726_c11_af83]
signal BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2726_c7_675a]
signal result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2726_c7_675a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2726_c7_675a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2726_c7_675a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2726_c7_675a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2732_c11_d60f]
signal BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2732_c7_92d9]
signal result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2732_c7_92d9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2732_c7_92d9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2732_c7_92d9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2736_c11_e46d]
signal BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2736_c7_9d77]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2736_c7_9d77]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_df93( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_value := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_stack_read := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_opc_done := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5
BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_left,
BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_right,
BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_return_output);

-- t8_MUX_uxn_opcodes_h_l2711_c2_e9a2
t8_MUX_uxn_opcodes_h_l2711_c2_e9a2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond,
t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue,
t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse,
t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2
result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond,
result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2
result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2
result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2
result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2
result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output);

-- printf_uxn_opcodes_h_l2712_c3_9a46_uxn_opcodes_h_l2712_c3_9a46
printf_uxn_opcodes_h_l2712_c3_9a46_uxn_opcodes_h_l2712_c3_9a46 : entity work.printf_uxn_opcodes_h_l2712_c3_9a46_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2712_c3_9a46_uxn_opcodes_h_l2712_c3_9a46_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c
BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_left,
BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_right,
BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output);

-- t8_MUX_uxn_opcodes_h_l2717_c7_e289
t8_MUX_uxn_opcodes_h_l2717_c7_e289 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2717_c7_e289_cond,
t8_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue,
t8_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse,
t8_MUX_uxn_opcodes_h_l2717_c7_e289_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289
result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_cond,
result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289
result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289
result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289
result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289
result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289
result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b
BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_left,
BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_right,
BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output);

-- t8_MUX_uxn_opcodes_h_l2720_c7_6f9b
t8_MUX_uxn_opcodes_h_l2720_c7_6f9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond,
t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue,
t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse,
t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b
result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond,
result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b
result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b
result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b
result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b
result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56
BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_left,
BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_right,
BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9
BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_left,
BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_right,
BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_return_output);

-- MUX_uxn_opcodes_h_l2724_c32_475a
MUX_uxn_opcodes_h_l2724_c32_475a : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2724_c32_475a_cond,
MUX_uxn_opcodes_h_l2724_c32_475a_iftrue,
MUX_uxn_opcodes_h_l2724_c32_475a_iffalse,
MUX_uxn_opcodes_h_l2724_c32_475a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83
BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_left,
BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_right,
BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a
result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_cond,
result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a
result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a
result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a
result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f
BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_left,
BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_right,
BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9
result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_cond,
result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9
result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9
result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d
BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_left,
BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_right,
BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77
result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77
result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_return_output,
 t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output,
 t8_MUX_uxn_opcodes_h_l2717_c7_e289_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output,
 t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_return_output,
 BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_return_output,
 MUX_uxn_opcodes_h_l2724_c32_475a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2714_c3_1d6a : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2712_c3_9a46_uxn_opcodes_h_l2712_c3_9a46_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2718_c3_6134 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2724_c32_475a_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2724_c32_475a_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2724_c32_475a_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2724_c32_475a_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2729_c3_6664 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2733_c3_9fd6 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2717_l2732_l2720_l2711_DUPLICATE_6284_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2717_l2711_l2726_DUPLICATE_affb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2717_l2720_l2711_DUPLICATE_8085_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2717_l2711_l2736_l2732_l2720_DUPLICATE_23cc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2717_l2720_DUPLICATE_296a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2717_l2736_l2732_l2726_l2720_DUPLICATE_89cc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2732_l2720_DUPLICATE_a6fa_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_df93_uxn_opcodes_h_l2707_l2741_DUPLICATE_5094_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2718_c3_6134 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2718_c3_6134;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_right := to_unsigned(4, 3);
     VAR_BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_right := to_unsigned(128, 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l2724_c32_475a_iftrue := signed(std_logic_vector(resize(to_unsigned(2, 2), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2733_c3_9fd6 := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2733_c3_9fd6;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2714_c3_1d6a := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2714_c3_1d6a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_right := to_unsigned(0, 1);
     VAR_BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_right := to_unsigned(0, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2729_c3_6664 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2729_c3_6664;
     VAR_MUX_uxn_opcodes_h_l2724_c32_475a_iffalse := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue := t8;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2717_l2732_l2720_l2711_DUPLICATE_6284 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2717_l2732_l2720_l2711_DUPLICATE_6284_return_output := result.stack_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2732_c11_d60f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2720_c11_557b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2711_c6_84f5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2717_l2720_DUPLICATE_296a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2717_l2720_DUPLICATE_296a_return_output := result.is_stack_read;

     -- BIN_OP_EQ[uxn_opcodes_h_l2726_c11_af83] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_left;
     BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_return_output := BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2717_c11_0f6c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l2724_c32_ef56] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_left;
     BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_return_output := BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2717_l2720_l2711_DUPLICATE_8085 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2717_l2720_l2711_DUPLICATE_8085_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2736_c11_e46d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2717_l2711_l2726_DUPLICATE_affb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2717_l2711_l2726_DUPLICATE_affb_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2732_l2720_DUPLICATE_a6fa LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2732_l2720_DUPLICATE_a6fa_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2717_l2711_l2736_l2732_l2720_DUPLICATE_23cc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2717_l2711_l2736_l2732_l2720_DUPLICATE_23cc_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2717_l2736_l2732_l2726_l2720_DUPLICATE_89cc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2717_l2736_l2732_l2726_l2720_DUPLICATE_89cc_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_left := VAR_BIN_OP_AND_uxn_opcodes_h_l2724_c32_ef56_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c6_84f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2717_c7_e289_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2717_c11_0f6c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2720_c11_557b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2726_c11_af83_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2732_c11_d60f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_e46d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2717_l2720_l2711_DUPLICATE_8085_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2717_l2720_l2711_DUPLICATE_8085_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2717_l2720_l2711_DUPLICATE_8085_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2717_l2736_l2732_l2726_l2720_DUPLICATE_89cc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2717_l2736_l2732_l2726_l2720_DUPLICATE_89cc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2717_l2736_l2732_l2726_l2720_DUPLICATE_89cc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2717_l2736_l2732_l2726_l2720_DUPLICATE_89cc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2717_l2736_l2732_l2726_l2720_DUPLICATE_89cc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2717_l2711_l2726_DUPLICATE_affb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2717_l2711_l2726_DUPLICATE_affb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2717_l2711_l2726_DUPLICATE_affb_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2717_l2720_DUPLICATE_296a_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2717_l2720_DUPLICATE_296a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2717_l2711_l2736_l2732_l2720_DUPLICATE_23cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2717_l2711_l2736_l2732_l2720_DUPLICATE_23cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2717_l2711_l2736_l2732_l2720_DUPLICATE_23cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2717_l2711_l2736_l2732_l2720_DUPLICATE_23cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2717_l2711_l2736_l2732_l2720_DUPLICATE_23cc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2732_l2720_DUPLICATE_a6fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2732_l2720_DUPLICATE_a6fa_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2717_l2732_l2720_l2711_DUPLICATE_6284_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2717_l2732_l2720_l2711_DUPLICATE_6284_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2717_l2732_l2720_l2711_DUPLICATE_6284_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2717_l2732_l2720_l2711_DUPLICATE_6284_return_output;
     -- result_stack_value_MUX[uxn_opcodes_h_l2732_c7_92d9] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output := result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l2724_c32_c2a9] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_left;
     BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_return_output := BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2720_c7_6f9b] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;

     -- t8_MUX[uxn_opcodes_h_l2720_c7_6f9b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond <= VAR_t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond;
     t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue;
     t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output := t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2711_c1_c79e] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2736_c7_9d77] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2736_c7_9d77] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2732_c7_92d9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2726_c7_675a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l2724_c32_475a_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l2724_c32_c2a9_return_output;
     VAR_printf_uxn_opcodes_h_l2712_c3_9a46_uxn_opcodes_h_l2712_c3_9a46_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2711_c1_c79e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2726_c7_675a_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_9d77_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2732_c7_92d9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output;

     -- printf_uxn_opcodes_h_l2712_c3_9a46[uxn_opcodes_h_l2712_c3_9a46] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2712_c3_9a46_uxn_opcodes_h_l2712_c3_9a46_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2712_c3_9a46_uxn_opcodes_h_l2712_c3_9a46_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2726_c7_675a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2726_c7_675a] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_return_output := result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2732_c7_92d9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output;

     -- t8_MUX[uxn_opcodes_h_l2717_c7_e289] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2717_c7_e289_cond <= VAR_t8_MUX_uxn_opcodes_h_l2717_c7_e289_cond;
     t8_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue;
     t8_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2717_c7_e289_return_output := t8_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;

     -- MUX[uxn_opcodes_h_l2724_c32_475a] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2724_c32_475a_cond <= VAR_MUX_uxn_opcodes_h_l2724_c32_475a_cond;
     MUX_uxn_opcodes_h_l2724_c32_475a_iftrue <= VAR_MUX_uxn_opcodes_h_l2724_c32_475a_iftrue;
     MUX_uxn_opcodes_h_l2724_c32_475a_iffalse <= VAR_MUX_uxn_opcodes_h_l2724_c32_475a_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2724_c32_475a_return_output := MUX_uxn_opcodes_h_l2724_c32_475a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2720_c7_6f9b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2717_c7_e289] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue := VAR_MUX_uxn_opcodes_h_l2724_c32_475a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2732_c7_92d9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2726_c7_675a_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2726_c7_675a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2717_c7_e289] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2711_c2_e9a2] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output;

     -- t8_MUX[uxn_opcodes_h_l2711_c2_e9a2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond <= VAR_t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond;
     t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue;
     t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output := t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2720_c7_6f9b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2726_c7_675a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2720_c7_6f9b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2720_c7_6f9b] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output := result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2726_c7_675a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2726_c7_675a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2726_c7_675a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2717_c7_e289] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2720_c7_6f9b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2711_c2_e9a2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2717_c7_e289] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2720_c7_6f9b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2717_c7_e289] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_return_output := result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2720_c7_6f9b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2717_c7_e289] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2711_c2_e9a2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2711_c2_e9a2] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output := result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2711_c2_e9a2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2717_c7_e289] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2717_c7_e289_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2711_c2_e9a2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2711_c2_e9a2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_df93_uxn_opcodes_h_l2707_l2741_DUPLICATE_5094 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_df93_uxn_opcodes_h_l2707_l2741_DUPLICATE_5094_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_df93(
     result,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c2_e9a2_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_df93_uxn_opcodes_h_l2707_l2741_DUPLICATE_5094_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_df93_uxn_opcodes_h_l2707_l2741_DUPLICATE_5094_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
