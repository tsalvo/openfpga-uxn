-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity gth_0CLK_441a128d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end gth_0CLK_441a128d;
architecture arch of gth_0CLK_441a128d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1809_c6_2494]
signal BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1809_c2_8f4d]
signal n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1809_c2_8f4d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1809_c2_8f4d]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1809_c2_8f4d]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1809_c2_8f4d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1809_c2_8f4d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1809_c2_8f4d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1809_c2_8f4d]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1809_c2_8f4d]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1809_c2_8f4d]
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1809_c2_8f4d]
signal t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1822_c11_acfd]
signal BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1822_c7_febd]
signal n8_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1822_c7_febd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1822_c7_febd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1822_c7_febd]
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1822_c7_febd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1822_c7_febd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1822_c7_febd]
signal t8_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1825_c11_1ea5]
signal BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1825_c7_94ae]
signal n8_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1825_c7_94ae]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1825_c7_94ae]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1825_c7_94ae]
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1825_c7_94ae]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1825_c7_94ae]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1825_c7_94ae]
signal t8_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1828_c11_30f2]
signal BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1828_c7_32fc]
signal n8_MUX_uxn_opcodes_h_l1828_c7_32fc_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1828_c7_32fc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1828_c7_32fc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1828_c7_32fc]
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1828_c7_32fc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1828_c7_32fc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1830_c30_a71f]
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_return_output : signed(3 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1833_c21_1ca0]
signal BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_right : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1833_c21_2d10]
signal MUX_uxn_opcodes_h_l1833_c21_2d10_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1833_c21_2d10_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1833_c21_2d10_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1833_c21_2d10_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8b52( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_left,
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_right,
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output);

-- n8_MUX_uxn_opcodes_h_l1809_c2_8f4d
n8_MUX_uxn_opcodes_h_l1809_c2_8f4d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond,
n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue,
n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse,
n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output);

-- t8_MUX_uxn_opcodes_h_l1809_c2_8f4d
t8_MUX_uxn_opcodes_h_l1809_c2_8f4d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond,
t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue,
t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse,
t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_left,
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_right,
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_return_output);

-- n8_MUX_uxn_opcodes_h_l1822_c7_febd
n8_MUX_uxn_opcodes_h_l1822_c7_febd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1822_c7_febd_cond,
n8_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue,
n8_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse,
n8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_cond,
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_return_output);

-- t8_MUX_uxn_opcodes_h_l1822_c7_febd
t8_MUX_uxn_opcodes_h_l1822_c7_febd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1822_c7_febd_cond,
t8_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue,
t8_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse,
t8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_left,
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_right,
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_return_output);

-- n8_MUX_uxn_opcodes_h_l1825_c7_94ae
n8_MUX_uxn_opcodes_h_l1825_c7_94ae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1825_c7_94ae_cond,
n8_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue,
n8_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse,
n8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_cond,
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output);

-- t8_MUX_uxn_opcodes_h_l1825_c7_94ae
t8_MUX_uxn_opcodes_h_l1825_c7_94ae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1825_c7_94ae_cond,
t8_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue,
t8_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse,
t8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_left,
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_right,
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_return_output);

-- n8_MUX_uxn_opcodes_h_l1828_c7_32fc
n8_MUX_uxn_opcodes_h_l1828_c7_32fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1828_c7_32fc_cond,
n8_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue,
n8_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse,
n8_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_cond,
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f
sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_ins,
sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_x,
sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_y,
sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0
BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0 : entity work.BIN_OP_GT_uint8_t_uint8_t_0CLK_380ecc95 port map (
BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_left,
BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_right,
BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_return_output);

-- MUX_uxn_opcodes_h_l1833_c21_2d10
MUX_uxn_opcodes_h_l1833_c21_2d10 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1833_c21_2d10_cond,
MUX_uxn_opcodes_h_l1833_c21_2d10_iftrue,
MUX_uxn_opcodes_h_l1833_c21_2d10_iffalse,
MUX_uxn_opcodes_h_l1833_c21_2d10_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output,
 n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
 t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_return_output,
 n8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_return_output,
 t8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_return_output,
 n8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output,
 t8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_return_output,
 n8_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output,
 sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_return_output,
 MUX_uxn_opcodes_h_l1833_c21_2d10_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1814_c3_60ee : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1819_c3_b15f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1823_c3_58d0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_febd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_94ae_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_32fc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1832_c3_bd9e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_2d10_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_2d10_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_2d10_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_2d10_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_53fb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_add5_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_6bc0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_418a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_9066_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l1837_l1805_DUPLICATE_7099_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_right := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1833_c21_2d10_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_y := resize(to_signed(-1, 2), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1819_c3_b15f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1819_c3_b15f;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1814_c3_60ee := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1814_c3_60ee;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_right := to_unsigned(2, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_right := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1833_c21_2d10_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1832_c3_bd9e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1832_c3_bd9e;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1823_c3_58d0 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1823_c3_58d0;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_418a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_418a_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1822_c11_acfd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_left;
     BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_return_output := BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1830_c30_a71f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_ins;
     sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_x;
     sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_return_output := sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1809_c2_8f4d_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_6bc0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_6bc0_return_output := result.is_stack_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1809_c2_8f4d_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1828_c11_30f2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_add5 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_add5_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1825_c11_1ea5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1809_c2_8f4d_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_9066 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_9066_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_53fb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_53fb_return_output := result.u8_value;

     -- BIN_OP_GT[uxn_opcodes_h_l1833_c21_1ca0] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_left;
     BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_return_output := BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1809_c2_8f4d_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1809_c6_2494] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_left;
     BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output := BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_2494_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_febd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_febd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_acfd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_94ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_94ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_1ea5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_32fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_30f2_return_output;
     VAR_MUX_uxn_opcodes_h_l1833_c21_2d10_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_1ca0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_add5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_add5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_add5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_418a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_418a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_418a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_6bc0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_6bc0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_6bc0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_9066_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_9066_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_53fb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_53fb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_53fb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_53fb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1809_c2_8f4d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1809_c2_8f4d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1809_c2_8f4d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1809_c2_8f4d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_a71f_return_output;
     -- n8_MUX[uxn_opcodes_h_l1828_c7_32fc] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1828_c7_32fc_cond <= VAR_n8_MUX_uxn_opcodes_h_l1828_c7_32fc_cond;
     n8_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue;
     n8_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output := n8_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1828_c7_32fc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output;

     -- MUX[uxn_opcodes_h_l1833_c21_2d10] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1833_c21_2d10_cond <= VAR_MUX_uxn_opcodes_h_l1833_c21_2d10_cond;
     MUX_uxn_opcodes_h_l1833_c21_2d10_iftrue <= VAR_MUX_uxn_opcodes_h_l1833_c21_2d10_iftrue;
     MUX_uxn_opcodes_h_l1833_c21_2d10_iffalse <= VAR_MUX_uxn_opcodes_h_l1833_c21_2d10_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1833_c21_2d10_return_output := MUX_uxn_opcodes_h_l1833_c21_2d10_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1828_c7_32fc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1828_c7_32fc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output;

     -- t8_MUX[uxn_opcodes_h_l1825_c7_94ae] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1825_c7_94ae_cond <= VAR_t8_MUX_uxn_opcodes_h_l1825_c7_94ae_cond;
     t8_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue;
     t8_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output := t8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1828_c7_32fc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue := VAR_MUX_uxn_opcodes_h_l1833_c21_2d10_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1825_c7_94ae] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;

     -- n8_MUX[uxn_opcodes_h_l1825_c7_94ae] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1825_c7_94ae_cond <= VAR_n8_MUX_uxn_opcodes_h_l1825_c7_94ae_cond;
     n8_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue;
     n8_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output := n8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1825_c7_94ae] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1825_c7_94ae] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1825_c7_94ae] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;

     -- t8_MUX[uxn_opcodes_h_l1822_c7_febd] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1822_c7_febd_cond <= VAR_t8_MUX_uxn_opcodes_h_l1822_c7_febd_cond;
     t8_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue;
     t8_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output := t8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1828_c7_32fc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output := result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_32fc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;
     -- t8_MUX[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond <= VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond;
     t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue;
     t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output := t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1825_c7_94ae] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output := result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1822_c7_febd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;

     -- n8_MUX[uxn_opcodes_h_l1822_c7_febd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1822_c7_febd_cond <= VAR_n8_MUX_uxn_opcodes_h_l1822_c7_febd_cond;
     n8_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue;
     n8_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output := n8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1822_c7_febd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1822_c7_febd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1822_c7_febd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_94ae_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output;
     -- n8_MUX[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond <= VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond;
     n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue;
     n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output := n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1822_c7_febd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_return_output := result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_febd_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1809_c2_8f4d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l1837_l1805_DUPLICATE_7099 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l1837_l1805_DUPLICATE_7099_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8b52(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_8f4d_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l1837_l1805_DUPLICATE_7099_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l1837_l1805_DUPLICATE_7099_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
