-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity mul_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end mul_0CLK_bacf6a1d;
architecture arch of mul_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1874_c6_1c62]
signal BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1874_c1_8dc8]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1874_c2_e391]
signal t8_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1874_c2_e391]
signal n8_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1874_c2_e391]
signal result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1874_c2_e391]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1874_c2_e391]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1874_c2_e391]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1874_c2_e391]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1874_c2_e391]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l1875_c3_e24f[uxn_opcodes_h_l1875_c3_e24f]
signal printf_uxn_opcodes_h_l1875_c3_e24f_uxn_opcodes_h_l1875_c3_e24f_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1879_c11_1276]
signal BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1879_c7_66a4]
signal t8_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1879_c7_66a4]
signal n8_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1879_c7_66a4]
signal result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1879_c7_66a4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1879_c7_66a4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1879_c7_66a4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1879_c7_66a4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1879_c7_66a4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1882_c11_c402]
signal BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1882_c7_b272]
signal t8_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1882_c7_b272]
signal n8_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1882_c7_b272]
signal result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1882_c7_b272]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1882_c7_b272]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1882_c7_b272]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1882_c7_b272]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1882_c7_b272]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1885_c11_305a]
signal BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1885_c7_8b50]
signal n8_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1885_c7_8b50]
signal result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1885_c7_8b50]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1885_c7_8b50]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1885_c7_8b50]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1885_c7_8b50]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1885_c7_8b50]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1888_c30_bd0e]
signal sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_return_output : signed(3 downto 0);

-- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1891_c21_49d2]
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_left : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_right : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1893_c11_e26f]
signal BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1893_c7_c651]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1893_c7_c651]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1893_c7_c651]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62
BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_left,
BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_right,
BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_return_output);

-- t8_MUX_uxn_opcodes_h_l1874_c2_e391
t8_MUX_uxn_opcodes_h_l1874_c2_e391 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1874_c2_e391_cond,
t8_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue,
t8_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse,
t8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output);

-- n8_MUX_uxn_opcodes_h_l1874_c2_e391
n8_MUX_uxn_opcodes_h_l1874_c2_e391 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1874_c2_e391_cond,
n8_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue,
n8_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse,
n8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391
result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_cond,
result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391
result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391
result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391
result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391
result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output);

-- printf_uxn_opcodes_h_l1875_c3_e24f_uxn_opcodes_h_l1875_c3_e24f
printf_uxn_opcodes_h_l1875_c3_e24f_uxn_opcodes_h_l1875_c3_e24f : entity work.printf_uxn_opcodes_h_l1875_c3_e24f_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1875_c3_e24f_uxn_opcodes_h_l1875_c3_e24f_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276
BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_left,
BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_right,
BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output);

-- t8_MUX_uxn_opcodes_h_l1879_c7_66a4
t8_MUX_uxn_opcodes_h_l1879_c7_66a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1879_c7_66a4_cond,
t8_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue,
t8_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse,
t8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output);

-- n8_MUX_uxn_opcodes_h_l1879_c7_66a4
n8_MUX_uxn_opcodes_h_l1879_c7_66a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1879_c7_66a4_cond,
n8_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue,
n8_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse,
n8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4
result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402
BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_left,
BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_right,
BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output);

-- t8_MUX_uxn_opcodes_h_l1882_c7_b272
t8_MUX_uxn_opcodes_h_l1882_c7_b272 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1882_c7_b272_cond,
t8_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue,
t8_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse,
t8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output);

-- n8_MUX_uxn_opcodes_h_l1882_c7_b272
n8_MUX_uxn_opcodes_h_l1882_c7_b272 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1882_c7_b272_cond,
n8_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue,
n8_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse,
n8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272
result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_cond,
result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272
result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272
result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272
result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272
result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a
BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_left,
BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_right,
BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_return_output);

-- n8_MUX_uxn_opcodes_h_l1885_c7_8b50
n8_MUX_uxn_opcodes_h_l1885_c7_8b50 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1885_c7_8b50_cond,
n8_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue,
n8_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse,
n8_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50
result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_cond,
result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50
result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e
sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_ins,
sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_x,
sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_y,
sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_return_output);

-- BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2 : entity work.BIN_OP_INFERRED_MULT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_left,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_right,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f
BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_left,
BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_right,
BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651
result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651
result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651
result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_return_output,
 t8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output,
 n8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output,
 t8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output,
 n8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output,
 t8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output,
 n8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_return_output,
 n8_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output,
 sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_return_output,
 BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1876_c3_4eff : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1875_c3_e24f_uxn_opcodes_h_l1875_c3_e24f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1880_c3_04cd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l1891_c3_7cac : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1890_c3_c203 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_dce5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_8271_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_44c0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_3d83_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1885_l1879_l1893_l1882_DUPLICATE_42a6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1885_l1882_DUPLICATE_314f_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1899_l1870_DUPLICATE_f0c6_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1876_c3_4eff := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1876_c3_4eff;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1880_c3_04cd := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1880_c3_04cd;
     VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1890_c3_c203 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1890_c3_c203;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_left := VAR_phase;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_dce5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_dce5_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1885_c11_305a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1874_c6_1c62] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_left;
     BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output := BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_3d83 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_3d83_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l1888_c30_bd0e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_ins;
     sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_x;
     sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_return_output := sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1893_c11_e26f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1879_c11_1276] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_left;
     BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output := BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_8271 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_8271_return_output := result.is_sp_shift;

     -- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1891_c21_49d2] LATENCY=0
     -- Inputs
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_left <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_left;
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_right <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_right;
     -- Outputs
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_return_output := BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1885_l1879_l1893_l1882_DUPLICATE_42a6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1885_l1879_l1893_l1882_DUPLICATE_42a6_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_44c0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_44c0_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1882_c11_c402] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_left;
     BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output := BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1885_l1882_DUPLICATE_314f LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1885_l1882_DUPLICATE_314f_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1874_c2_e391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1874_c2_e391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_1c62_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1879_c7_66a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1879_c7_66a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_1276_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1882_c7_b272_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1882_c7_b272_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_c402_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1885_c7_8b50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_305a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_e26f_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l1891_c3_7cac := resize(VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_49d2_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_3d83_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_3d83_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_3d83_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_3d83_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1885_l1879_l1893_l1882_DUPLICATE_42a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1885_l1879_l1893_l1882_DUPLICATE_42a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1885_l1879_l1893_l1882_DUPLICATE_42a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1885_l1879_l1893_l1882_DUPLICATE_42a6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_8271_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_8271_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_8271_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_8271_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_44c0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_44c0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_44c0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1874_l1879_l1893_l1882_DUPLICATE_44c0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1885_l1882_DUPLICATE_314f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1885_l1882_DUPLICATE_314f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_dce5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_dce5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_dce5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1874_l1885_l1879_l1882_DUPLICATE_dce5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_bd0e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue := VAR_result_u8_value_uxn_opcodes_h_l1891_c3_7cac;
     -- result_u8_value_MUX[uxn_opcodes_h_l1885_c7_8b50] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output := result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;

     -- n8_MUX[uxn_opcodes_h_l1885_c7_8b50] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1885_c7_8b50_cond <= VAR_n8_MUX_uxn_opcodes_h_l1885_c7_8b50_cond;
     n8_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue;
     n8_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output := n8_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1885_c7_8b50] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1885_c7_8b50] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1893_c7_c651] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1893_c7_c651] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1893_c7_c651] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1874_c1_8dc8] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_return_output;

     -- t8_MUX[uxn_opcodes_h_l1882_c7_b272] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1882_c7_b272_cond <= VAR_t8_MUX_uxn_opcodes_h_l1882_c7_b272_cond;
     t8_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue;
     t8_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output := t8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l1875_c3_e24f_uxn_opcodes_h_l1875_c3_e24f_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_8dc8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c651_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c651_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c651_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1885_c7_8b50] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;

     -- t8_MUX[uxn_opcodes_h_l1879_c7_66a4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1879_c7_66a4_cond <= VAR_t8_MUX_uxn_opcodes_h_l1879_c7_66a4_cond;
     t8_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue;
     t8_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output := t8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1882_c7_b272] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_return_output := result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1882_c7_b272] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1885_c7_8b50] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;

     -- printf_uxn_opcodes_h_l1875_c3_e24f[uxn_opcodes_h_l1875_c3_e24f] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1875_c3_e24f_uxn_opcodes_h_l1875_c3_e24f_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1875_c3_e24f_uxn_opcodes_h_l1875_c3_e24f_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- n8_MUX[uxn_opcodes_h_l1882_c7_b272] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1882_c7_b272_cond <= VAR_n8_MUX_uxn_opcodes_h_l1882_c7_b272_cond;
     n8_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue;
     n8_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output := n8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1885_c7_8b50] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1882_c7_b272] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_8b50_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1879_c7_66a4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1879_c7_66a4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;

     -- t8_MUX[uxn_opcodes_h_l1874_c2_e391] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1874_c2_e391_cond <= VAR_t8_MUX_uxn_opcodes_h_l1874_c2_e391_cond;
     t8_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue;
     t8_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output := t8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1879_c7_66a4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1882_c7_b272] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;

     -- n8_MUX[uxn_opcodes_h_l1879_c7_66a4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1879_c7_66a4_cond <= VAR_n8_MUX_uxn_opcodes_h_l1879_c7_66a4_cond;
     n8_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue;
     n8_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output := n8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1882_c7_b272] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1882_c7_b272] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_b272_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1874_c2_e391] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1879_c7_66a4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1879_c7_66a4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1879_c7_66a4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1874_c2_e391] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1874_c2_e391_cond <= VAR_n8_MUX_uxn_opcodes_h_l1874_c2_e391_cond;
     n8_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue;
     n8_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output := n8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1874_c2_e391] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1874_c2_e391] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_return_output := result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1874_c2_e391_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_66a4_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1874_c2_e391] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1874_c2_e391] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1874_c2_e391] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1899_l1870_DUPLICATE_f0c6 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1899_l1870_DUPLICATE_f0c6_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_e391_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_e391_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_e391_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_e391_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_e391_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1899_l1870_DUPLICATE_f0c6_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1899_l1870_DUPLICATE_f0c6_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
