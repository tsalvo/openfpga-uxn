-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity and_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end and_0CLK_bacf6a1d;
architecture arch of and_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l869_c6_5c68]
signal BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l869_c1_7b1d]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l869_c2_872c]
signal n8_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l869_c2_872c]
signal t8_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l869_c2_872c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l869_c2_872c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l869_c2_872c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l869_c2_872c]
signal result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l869_c2_872c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l869_c2_872c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l870_c3_c40e[uxn_opcodes_h_l870_c3_c40e]
signal printf_uxn_opcodes_h_l870_c3_c40e_uxn_opcodes_h_l870_c3_c40e_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l874_c11_3d32]
signal BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l874_c7_faf0]
signal n8_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l874_c7_faf0]
signal t8_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l874_c7_faf0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l874_c7_faf0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l874_c7_faf0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l874_c7_faf0]
signal result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l874_c7_faf0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l874_c7_faf0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l877_c11_2b87]
signal BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l877_c7_cb97]
signal n8_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l877_c7_cb97]
signal t8_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l877_c7_cb97]
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l877_c7_cb97]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l877_c7_cb97]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l877_c7_cb97]
signal result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l877_c7_cb97]
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l877_c7_cb97]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l880_c11_d129]
signal BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l880_c7_c191]
signal n8_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l880_c7_c191_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l880_c7_c191]
signal result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l880_c7_c191]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l880_c7_c191]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l880_c7_c191]
signal result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l880_c7_c191]
signal result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l880_c7_c191]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l883_c30_9bae]
signal sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_return_output : signed(3 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l886_c21_1043]
signal BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l888_c11_df5b]
signal BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l888_c7_36b3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l888_c7_36b3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l888_c7_36b3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c551( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68
BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_left,
BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_right,
BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_return_output);

-- n8_MUX_uxn_opcodes_h_l869_c2_872c
n8_MUX_uxn_opcodes_h_l869_c2_872c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l869_c2_872c_cond,
n8_MUX_uxn_opcodes_h_l869_c2_872c_iftrue,
n8_MUX_uxn_opcodes_h_l869_c2_872c_iffalse,
n8_MUX_uxn_opcodes_h_l869_c2_872c_return_output);

-- t8_MUX_uxn_opcodes_h_l869_c2_872c
t8_MUX_uxn_opcodes_h_l869_c2_872c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l869_c2_872c_cond,
t8_MUX_uxn_opcodes_h_l869_c2_872c_iftrue,
t8_MUX_uxn_opcodes_h_l869_c2_872c_iffalse,
t8_MUX_uxn_opcodes_h_l869_c2_872c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c
result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c
result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_cond,
result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c
result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output);

-- printf_uxn_opcodes_h_l870_c3_c40e_uxn_opcodes_h_l870_c3_c40e
printf_uxn_opcodes_h_l870_c3_c40e_uxn_opcodes_h_l870_c3_c40e : entity work.printf_uxn_opcodes_h_l870_c3_c40e_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l870_c3_c40e_uxn_opcodes_h_l870_c3_c40e_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32
BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_left,
BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_right,
BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output);

-- n8_MUX_uxn_opcodes_h_l874_c7_faf0
n8_MUX_uxn_opcodes_h_l874_c7_faf0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l874_c7_faf0_cond,
n8_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue,
n8_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse,
n8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output);

-- t8_MUX_uxn_opcodes_h_l874_c7_faf0
t8_MUX_uxn_opcodes_h_l874_c7_faf0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l874_c7_faf0_cond,
t8_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue,
t8_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse,
t8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0
result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0
result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0
result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_cond,
result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0
result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0
result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87
BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_left,
BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_right,
BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output);

-- n8_MUX_uxn_opcodes_h_l877_c7_cb97
n8_MUX_uxn_opcodes_h_l877_c7_cb97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l877_c7_cb97_cond,
n8_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue,
n8_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse,
n8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output);

-- t8_MUX_uxn_opcodes_h_l877_c7_cb97
t8_MUX_uxn_opcodes_h_l877_c7_cb97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l877_c7_cb97_cond,
t8_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue,
t8_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse,
t8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97
result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_cond,
result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129
BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_left,
BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_right,
BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_return_output);

-- n8_MUX_uxn_opcodes_h_l880_c7_c191
n8_MUX_uxn_opcodes_h_l880_c7_c191 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l880_c7_c191_cond,
n8_MUX_uxn_opcodes_h_l880_c7_c191_iftrue,
n8_MUX_uxn_opcodes_h_l880_c7_c191_iffalse,
n8_MUX_uxn_opcodes_h_l880_c7_c191_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191
result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191
result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191
result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_cond,
result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191
result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191
result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output);

-- sp_relative_shift_uxn_opcodes_h_l883_c30_9bae
sp_relative_shift_uxn_opcodes_h_l883_c30_9bae : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_ins,
sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_x,
sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_y,
sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l886_c21_1043
BIN_OP_AND_uxn_opcodes_h_l886_c21_1043 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_left,
BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_right,
BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b
BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_left,
BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_right,
BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_return_output,
 n8_MUX_uxn_opcodes_h_l869_c2_872c_return_output,
 t8_MUX_uxn_opcodes_h_l869_c2_872c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output,
 n8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output,
 t8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output,
 n8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output,
 t8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_return_output,
 n8_MUX_uxn_opcodes_h_l880_c7_c191_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output,
 sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_return_output,
 BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l871_c3_e5e9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l870_c3_c40e_uxn_opcodes_h_l870_c3_c40e_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l875_c3_65e0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l880_c7_c191_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l885_c3_0ca4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_e529_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_1551_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_617e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_eeb8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l874_l888_l877_l880_DUPLICATE_ada5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l877_l880_DUPLICATE_bc03_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l865_l894_DUPLICATE_4980_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l871_c3_e5e9 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l871_c3_e5e9;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_right := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l875_c3_65e0 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l875_c3_65e0;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l885_c3_0ca4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l885_c3_0ca4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l869_c2_872c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l880_c7_c191_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_left := VAR_phase;
     VAR_BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l880_c7_c191_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l869_c2_872c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l888_c11_df5b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_left;
     BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_return_output := BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_617e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_617e_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_eeb8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_eeb8_return_output := result.is_sp_shift;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_1551 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_1551_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_e529 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_e529_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l874_c11_3d32] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_left;
     BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output := BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l883_c30_9bae] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_ins;
     sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_x <= VAR_sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_x;
     sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_y <= VAR_sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_return_output := sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l877_c11_2b87] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_left;
     BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output := BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l880_c11_d129] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_left;
     BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_return_output := BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l886_c21_1043] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_left;
     BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_return_output := BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l869_c6_5c68] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_left;
     BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output := BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l874_l888_l877_l880_DUPLICATE_ada5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l874_l888_l877_l880_DUPLICATE_ada5_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l877_l880_DUPLICATE_bc03 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l877_l880_DUPLICATE_bc03_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_iftrue := VAR_BIN_OP_AND_uxn_opcodes_h_l886_c21_1043_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l869_c2_872c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l869_c2_872c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c6_5c68_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l874_c7_faf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l874_c7_faf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_3d32_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l877_c7_cb97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l877_c7_cb97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_2b87_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l880_c7_c191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_d129_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_df5b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_1551_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_1551_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_1551_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_1551_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l874_l888_l877_l880_DUPLICATE_ada5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l874_l888_l877_l880_DUPLICATE_ada5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l874_l888_l877_l880_DUPLICATE_ada5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l874_l888_l877_l880_DUPLICATE_ada5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_eeb8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_eeb8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_eeb8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_eeb8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_e529_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_e529_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_e529_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l874_l888_l877_l869_DUPLICATE_e529_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l877_l880_DUPLICATE_bc03_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l877_l880_DUPLICATE_bc03_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_617e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_617e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_617e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l874_l877_l869_l880_DUPLICATE_617e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l883_c30_9bae_return_output;
     -- t8_MUX[uxn_opcodes_h_l877_c7_cb97] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l877_c7_cb97_cond <= VAR_t8_MUX_uxn_opcodes_h_l877_c7_cb97_cond;
     t8_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue;
     t8_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output := t8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l888_c7_36b3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_return_output;

     -- n8_MUX[uxn_opcodes_h_l880_c7_c191] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l880_c7_c191_cond <= VAR_n8_MUX_uxn_opcodes_h_l880_c7_c191_cond;
     n8_MUX_uxn_opcodes_h_l880_c7_c191_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l880_c7_c191_iftrue;
     n8_MUX_uxn_opcodes_h_l880_c7_c191_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l880_c7_c191_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l880_c7_c191_return_output := n8_MUX_uxn_opcodes_h_l880_c7_c191_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l880_c7_c191] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l869_c1_7b1d] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l888_c7_36b3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l880_c7_c191] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l888_c7_36b3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l880_c7_c191] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_cond;
     result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_return_output := result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l870_c3_c40e_uxn_opcodes_h_l870_c3_c40e_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l869_c1_7b1d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse := VAR_n8_MUX_uxn_opcodes_h_l880_c7_c191_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_36b3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_36b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_36b3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l880_c7_c191_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l880_c7_c191_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l880_c7_c191] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l880_c7_c191] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_return_output;

     -- printf_uxn_opcodes_h_l870_c3_c40e[uxn_opcodes_h_l870_c3_c40e] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l870_c3_c40e_uxn_opcodes_h_l870_c3_c40e_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l870_c3_c40e_uxn_opcodes_h_l870_c3_c40e_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- t8_MUX[uxn_opcodes_h_l874_c7_faf0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l874_c7_faf0_cond <= VAR_t8_MUX_uxn_opcodes_h_l874_c7_faf0_cond;
     t8_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue;
     t8_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output := t8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;

     -- n8_MUX[uxn_opcodes_h_l877_c7_cb97] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l877_c7_cb97_cond <= VAR_n8_MUX_uxn_opcodes_h_l877_c7_cb97_cond;
     n8_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue;
     n8_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output := n8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l877_c7_cb97] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l877_c7_cb97] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l880_c7_c191] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l877_c7_cb97] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_cond;
     result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_return_output := result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_c191_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_c191_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_c191_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l869_c2_872c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l877_c7_cb97] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l877_c7_cb97] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;

     -- t8_MUX[uxn_opcodes_h_l869_c2_872c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l869_c2_872c_cond <= VAR_t8_MUX_uxn_opcodes_h_l869_c2_872c_cond;
     t8_MUX_uxn_opcodes_h_l869_c2_872c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l869_c2_872c_iftrue;
     t8_MUX_uxn_opcodes_h_l869_c2_872c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l869_c2_872c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l869_c2_872c_return_output := t8_MUX_uxn_opcodes_h_l869_c2_872c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l874_c7_faf0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l874_c7_faf0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;

     -- n8_MUX[uxn_opcodes_h_l874_c7_faf0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l874_c7_faf0_cond <= VAR_n8_MUX_uxn_opcodes_h_l874_c7_faf0_cond;
     n8_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue;
     n8_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output := n8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l874_c7_faf0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_return_output := result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l877_c7_cb97] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l869_c2_872c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_cb97_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l869_c2_872c_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l869_c2_872c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_return_output := result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l869_c2_872c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l874_c7_faf0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l874_c7_faf0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l869_c2_872c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_return_output;

     -- n8_MUX[uxn_opcodes_h_l869_c2_872c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l869_c2_872c_cond <= VAR_n8_MUX_uxn_opcodes_h_l869_c2_872c_cond;
     n8_MUX_uxn_opcodes_h_l869_c2_872c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l869_c2_872c_iftrue;
     n8_MUX_uxn_opcodes_h_l869_c2_872c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l869_c2_872c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l869_c2_872c_return_output := n8_MUX_uxn_opcodes_h_l869_c2_872c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l874_c7_faf0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l869_c2_872c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_faf0_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l869_c2_872c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l869_c2_872c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l869_c2_872c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l865_l894_DUPLICATE_4980 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l865_l894_DUPLICATE_4980_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c551(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c2_872c_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c2_872c_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c2_872c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c2_872c_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c2_872c_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l865_l894_DUPLICATE_4980_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l865_l894_DUPLICATE_4980_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
