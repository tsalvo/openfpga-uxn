-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity sth_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth_0CLK_85d5529e;
architecture arch of sth_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2259_c6_40a5]
signal BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2259_c1_94dd]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2259_c2_6e90]
signal t8_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2259_c2_6e90]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2259_c2_6e90]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2259_c2_6e90]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2259_c2_6e90]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2259_c2_6e90]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2259_c2_6e90]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2259_c2_6e90]
signal result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2260_c3_f7b6[uxn_opcodes_h_l2260_c3_f7b6]
signal printf_uxn_opcodes_h_l2260_c3_f7b6_uxn_opcodes_h_l2260_c3_f7b6_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2264_c11_e9a7]
signal BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2264_c7_d8a8]
signal t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2264_c7_d8a8]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2264_c7_d8a8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2264_c7_d8a8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2264_c7_d8a8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2264_c7_d8a8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2264_c7_d8a8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2264_c7_d8a8]
signal result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2267_c11_5ad8]
signal BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2267_c7_2b48]
signal t8_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2267_c7_2b48]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2267_c7_2b48]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2267_c7_2b48]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2267_c7_2b48]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2267_c7_2b48]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2267_c7_2b48]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2267_c7_2b48]
signal result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2270_c30_ad38]
signal sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2272_c11_d5d6]
signal BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2272_c7_b72b]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2272_c7_b72b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2272_c7_b72b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2272_c7_b72b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2272_c7_b72b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2272_c7_b72b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2272_c7_b72b]
signal result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2279_c11_86ea]
signal BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2279_c7_2cca]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2279_c7_2cca]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2279_c7_2cca]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2279_c7_2cca]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_10dd( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_index_flipped := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.u8_value := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5
BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_left,
BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_right,
BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_return_output);

-- t8_MUX_uxn_opcodes_h_l2259_c2_6e90
t8_MUX_uxn_opcodes_h_l2259_c2_6e90 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2259_c2_6e90_cond,
t8_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue,
t8_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse,
t8_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90
result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_cond,
result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output);

-- printf_uxn_opcodes_h_l2260_c3_f7b6_uxn_opcodes_h_l2260_c3_f7b6
printf_uxn_opcodes_h_l2260_c3_f7b6_uxn_opcodes_h_l2260_c3_f7b6 : entity work.printf_uxn_opcodes_h_l2260_c3_f7b6_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2260_c3_f7b6_uxn_opcodes_h_l2260_c3_f7b6_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7
BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_left,
BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_right,
BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output);

-- t8_MUX_uxn_opcodes_h_l2264_c7_d8a8
t8_MUX_uxn_opcodes_h_l2264_c7_d8a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond,
t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue,
t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse,
t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8
result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8
BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_left,
BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_right,
BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output);

-- t8_MUX_uxn_opcodes_h_l2267_c7_2b48
t8_MUX_uxn_opcodes_h_l2267_c7_2b48 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2267_c7_2b48_cond,
t8_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue,
t8_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse,
t8_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48
result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48
result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48
result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48
result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48
result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_cond,
result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38
sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_ins,
sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_x,
sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_y,
sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6
BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_left,
BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_right,
BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b
result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b
result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea
BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_left,
BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_right,
BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca
result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca
result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca
result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_return_output,
 t8_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output,
 t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output,
 t8_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output,
 sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2261_c3_bd71 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2260_c3_f7b6_uxn_opcodes_h_l2260_c3_f7b6_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2265_c3_0d8b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2276_c3_9a05 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2274_c3_e830 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_8da5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_54a2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2264_l2279_l2259_l2272_DUPLICATE_4cd1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2264_l2259_l2272_DUPLICATE_fb43_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2264_l2267_l2259_l2272_DUPLICATE_069f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2272_DUPLICATE_bb56_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2267_l2272_DUPLICATE_10c4_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_10dd_uxn_opcodes_h_l2255_l2286_DUPLICATE_c289_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2261_c3_bd71 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2261_c3_bd71;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2274_c3_e830 := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2274_c3_e830;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2276_c3_9a05 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2276_c3_9a05;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2265_c3_0d8b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2265_c3_0d8b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_right := to_unsigned(3, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse := t8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2267_l2272_DUPLICATE_10c4 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2267_l2272_DUPLICATE_10c4_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2279_c11_86ea] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_left;
     BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_return_output := BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2267_c11_5ad8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2264_l2267_l2259_l2272_DUPLICATE_069f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2264_l2267_l2259_l2272_DUPLICATE_069f_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_8da5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_8da5_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2272_DUPLICATE_bb56 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2272_DUPLICATE_bb56_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2272_c11_d5d6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_54a2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_54a2_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l2270_c30_ad38] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_ins;
     sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_x;
     sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_return_output := sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2259_c6_40a5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2264_c11_e9a7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_left;
     BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output := BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2264_l2259_l2272_DUPLICATE_fb43 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2264_l2259_l2272_DUPLICATE_fb43_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2264_l2279_l2259_l2272_DUPLICATE_4cd1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2264_l2279_l2259_l2272_DUPLICATE_4cd1_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2259_c2_6e90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2259_c6_40a5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2264_c11_e9a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2267_c7_2b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2267_c11_5ad8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2272_c11_d5d6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2279_c11_86ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2264_l2259_l2272_DUPLICATE_fb43_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2264_l2259_l2272_DUPLICATE_fb43_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2264_l2259_l2272_DUPLICATE_fb43_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2272_DUPLICATE_bb56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2272_DUPLICATE_bb56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2272_DUPLICATE_bb56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2272_DUPLICATE_bb56_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2264_l2279_l2259_l2272_DUPLICATE_4cd1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2264_l2279_l2259_l2272_DUPLICATE_4cd1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2264_l2279_l2259_l2272_DUPLICATE_4cd1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2264_l2279_l2259_l2272_DUPLICATE_4cd1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_8da5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_8da5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_8da5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_8da5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_54a2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_54a2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_54a2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2264_l2279_l2267_l2259_DUPLICATE_54a2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2267_l2272_DUPLICATE_10c4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2267_l2272_DUPLICATE_10c4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2264_l2267_l2259_l2272_DUPLICATE_069f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2264_l2267_l2259_l2272_DUPLICATE_069f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2264_l2267_l2259_l2272_DUPLICATE_069f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2264_l2267_l2259_l2272_DUPLICATE_069f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2270_c30_ad38_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2279_c7_2cca] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2272_c7_b72b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;

     -- t8_MUX[uxn_opcodes_h_l2267_c7_2b48] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2267_c7_2b48_cond <= VAR_t8_MUX_uxn_opcodes_h_l2267_c7_2b48_cond;
     t8_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue;
     t8_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output := t8_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2272_c7_b72b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2279_c7_2cca] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2259_c1_94dd] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2272_c7_b72b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2279_c7_2cca] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2279_c7_2cca] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2260_c3_f7b6_uxn_opcodes_h_l2260_c3_f7b6_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2259_c1_94dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2279_c7_2cca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2272_c7_b72b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2272_c7_b72b] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2272_c7_b72b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2272_c7_b72b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2267_c7_2b48] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;

     -- t8_MUX[uxn_opcodes_h_l2264_c7_d8a8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond <= VAR_t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond;
     t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue;
     t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output := t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;

     -- printf_uxn_opcodes_h_l2260_c3_f7b6[uxn_opcodes_h_l2260_c3_f7b6] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2260_c3_f7b6_uxn_opcodes_h_l2260_c3_f7b6_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2260_c3_f7b6_uxn_opcodes_h_l2260_c3_f7b6_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2267_c7_2b48] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2267_c7_2b48] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output := result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2272_c7_b72b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2264_c7_d8a8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2264_c7_d8a8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;

     -- t8_MUX[uxn_opcodes_h_l2259_c2_6e90] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2259_c2_6e90_cond <= VAR_t8_MUX_uxn_opcodes_h_l2259_c2_6e90_cond;
     t8_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue;
     t8_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output := t8_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2267_c7_2b48] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2264_c7_d8a8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2267_c7_2b48] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2267_c7_2b48] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2267_c7_2b48] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2267_c7_2b48_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2259_c2_6e90] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2259_c2_6e90] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output := result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2259_c2_6e90] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2264_c7_d8a8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2264_c7_d8a8] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2264_c7_d8a8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2264_c7_d8a8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2264_c7_d8a8_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2259_c2_6e90] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2259_c2_6e90] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2259_c2_6e90] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2259_c2_6e90] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_10dd_uxn_opcodes_h_l2255_l2286_DUPLICATE_c289 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_10dd_uxn_opcodes_h_l2255_l2286_DUPLICATE_c289_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_10dd(
     result,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2259_c2_6e90_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_10dd_uxn_opcodes_h_l2255_l2286_DUPLICATE_c289_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_10dd_uxn_opcodes_h_l2255_l2286_DUPLICATE_c289_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
