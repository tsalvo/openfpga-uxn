-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity gth_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end gth_0CLK_226c8821;
architecture arch of gth_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1809_c6_4ddd]
signal BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1809_c2_bab7]
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1809_c2_bab7]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1809_c2_bab7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1809_c2_bab7]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1809_c2_bab7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1809_c2_bab7]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1809_c2_bab7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1809_c2_bab7]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1809_c2_bab7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1809_c2_bab7]
signal n8_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1809_c2_bab7]
signal t8_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1822_c11_5878]
signal BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1822_c7_d6d6]
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1822_c7_d6d6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1822_c7_d6d6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1822_c7_d6d6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1822_c7_d6d6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1822_c7_d6d6]
signal n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1822_c7_d6d6]
signal t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1825_c11_8890]
signal BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1825_c7_f7c3]
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1825_c7_f7c3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1825_c7_f7c3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1825_c7_f7c3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1825_c7_f7c3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1825_c7_f7c3]
signal n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1825_c7_f7c3]
signal t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1828_c11_f0b7]
signal BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1828_c7_9124]
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1828_c7_9124]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1828_c7_9124]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1828_c7_9124]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1828_c7_9124]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1828_c7_9124]
signal n8_MUX_uxn_opcodes_h_l1828_c7_9124_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1828_c7_9124_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1830_c30_b044]
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_return_output : signed(3 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1833_c21_e65c]
signal BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_right : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1833_c21_7b51]
signal MUX_uxn_opcodes_h_l1833_c21_7b51_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1833_c21_7b51_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1833_c21_7b51_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1833_c21_7b51_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_922a( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_pc_updated := ref_toks_6;
      base.is_opc_done := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_left,
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_right,
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_cond,
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output);

-- n8_MUX_uxn_opcodes_h_l1809_c2_bab7
n8_MUX_uxn_opcodes_h_l1809_c2_bab7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1809_c2_bab7_cond,
n8_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue,
n8_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse,
n8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output);

-- t8_MUX_uxn_opcodes_h_l1809_c2_bab7
t8_MUX_uxn_opcodes_h_l1809_c2_bab7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1809_c2_bab7_cond,
t8_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue,
t8_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse,
t8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_left,
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_right,
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond,
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output);

-- n8_MUX_uxn_opcodes_h_l1822_c7_d6d6
n8_MUX_uxn_opcodes_h_l1822_c7_d6d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond,
n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue,
n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse,
n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output);

-- t8_MUX_uxn_opcodes_h_l1822_c7_d6d6
t8_MUX_uxn_opcodes_h_l1822_c7_d6d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond,
t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue,
t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse,
t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_left,
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_right,
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond,
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output);

-- n8_MUX_uxn_opcodes_h_l1825_c7_f7c3
n8_MUX_uxn_opcodes_h_l1825_c7_f7c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond,
n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue,
n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse,
n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output);

-- t8_MUX_uxn_opcodes_h_l1825_c7_f7c3
t8_MUX_uxn_opcodes_h_l1825_c7_f7c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond,
t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue,
t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse,
t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_left,
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_right,
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_cond,
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_return_output);

-- n8_MUX_uxn_opcodes_h_l1828_c7_9124
n8_MUX_uxn_opcodes_h_l1828_c7_9124 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1828_c7_9124_cond,
n8_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue,
n8_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse,
n8_MUX_uxn_opcodes_h_l1828_c7_9124_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1830_c30_b044
sp_relative_shift_uxn_opcodes_h_l1830_c30_b044 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_ins,
sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_x,
sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_y,
sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c
BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c : entity work.BIN_OP_GT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_left,
BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_right,
BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_return_output);

-- MUX_uxn_opcodes_h_l1833_c21_7b51
MUX_uxn_opcodes_h_l1833_c21_7b51 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1833_c21_7b51_cond,
MUX_uxn_opcodes_h_l1833_c21_7b51_iftrue,
MUX_uxn_opcodes_h_l1833_c21_7b51_iffalse,
MUX_uxn_opcodes_h_l1833_c21_7b51_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
 n8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
 t8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output,
 n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output,
 t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output,
 n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output,
 t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_return_output,
 n8_MUX_uxn_opcodes_h_l1828_c7_9124_return_output,
 sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_return_output,
 MUX_uxn_opcodes_h_l1833_c21_7b51_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1819_c3_1c60 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1814_c3_ce41 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_bab7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1823_c3_5caa : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_9124_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1832_c3_af57 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_9124_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_7b51_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_7b51_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_7b51_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_7b51_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1828_l1822_l1825_DUPLICATE_5784_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_0af3_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_b3fe_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_732d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1828_l1825_DUPLICATE_01e2_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1837_l1805_DUPLICATE_6ea5_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1814_c3_ce41 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1814_c3_ce41;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1832_c3_af57 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1832_c3_af57;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1833_c21_7b51_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1819_c3_1c60 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1819_c3_1c60;
     VAR_MUX_uxn_opcodes_h_l1833_c21_7b51_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1823_c3_5caa := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1823_c3_5caa;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1825_c11_8890] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_left;
     BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_return_output := BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1809_c2_bab7_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_732d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_732d_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1828_l1825_DUPLICATE_01e2 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1828_l1825_DUPLICATE_01e2_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l1830_c30_b044] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_ins;
     sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_x;
     sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_return_output := sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_0af3 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_0af3_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1828_c11_f0b7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_left;
     BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_return_output := BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1828_l1822_l1825_DUPLICATE_5784 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1828_l1822_l1825_DUPLICATE_5784_return_output := result.u8_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1809_c2_bab7_return_output := result.is_ram_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1809_c2_bab7_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1822_c11_5878] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_left;
     BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_return_output := BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1809_c6_4ddd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_left;
     BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output := BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1809_c2_bab7_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_b3fe LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_b3fe_return_output := result.is_opc_done;

     -- BIN_OP_GT[uxn_opcodes_h_l1833_c21_e65c] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_left;
     BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_return_output := BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_bab7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_bab7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_4ddd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_5878_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_8890_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_9124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_f0b7_return_output;
     VAR_MUX_uxn_opcodes_h_l1833_c21_7b51_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_e65c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_0af3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_0af3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_0af3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_b3fe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_b3fe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_b3fe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_732d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_732d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1828_l1822_l1825_DUPLICATE_732d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1828_l1825_DUPLICATE_01e2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1828_l1825_DUPLICATE_01e2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1828_l1822_l1825_DUPLICATE_5784_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1828_l1822_l1825_DUPLICATE_5784_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1828_l1822_l1825_DUPLICATE_5784_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1809_l1828_l1822_l1825_DUPLICATE_5784_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1809_c2_bab7_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1809_c2_bab7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1809_c2_bab7_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1809_c2_bab7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_b044_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1828_c7_9124] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1828_c7_9124] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1828_c7_9124] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1828_c7_9124] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_return_output;

     -- n8_MUX[uxn_opcodes_h_l1828_c7_9124] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1828_c7_9124_cond <= VAR_n8_MUX_uxn_opcodes_h_l1828_c7_9124_cond;
     n8_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue;
     n8_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_9124_return_output := n8_MUX_uxn_opcodes_h_l1828_c7_9124_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output;

     -- t8_MUX[uxn_opcodes_h_l1825_c7_f7c3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond <= VAR_t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond;
     t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue;
     t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output := t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output;

     -- MUX[uxn_opcodes_h_l1833_c21_7b51] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1833_c21_7b51_cond <= VAR_MUX_uxn_opcodes_h_l1833_c21_7b51_cond;
     MUX_uxn_opcodes_h_l1833_c21_7b51_iftrue <= VAR_MUX_uxn_opcodes_h_l1833_c21_7b51_iftrue;
     MUX_uxn_opcodes_h_l1833_c21_7b51_iffalse <= VAR_MUX_uxn_opcodes_h_l1833_c21_7b51_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1833_c21_7b51_return_output := MUX_uxn_opcodes_h_l1833_c21_7b51_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue := VAR_MUX_uxn_opcodes_h_l1833_c21_7b51_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1828_c7_9124_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_9124_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_9124_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_9124_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_9124_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1825_c7_f7c3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;

     -- n8_MUX[uxn_opcodes_h_l1825_c7_f7c3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond <= VAR_n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond;
     n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue;
     n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output := n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1828_c7_9124] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_return_output := result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1825_c7_f7c3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1825_c7_f7c3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;

     -- t8_MUX[uxn_opcodes_h_l1822_c7_d6d6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond <= VAR_t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond;
     t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue;
     t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output := t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1825_c7_f7c3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_9124_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1822_c7_d6d6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1822_c7_d6d6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;

     -- n8_MUX[uxn_opcodes_h_l1822_c7_d6d6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond <= VAR_n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond;
     n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue;
     n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output := n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1822_c7_d6d6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;

     -- t8_MUX[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1809_c2_bab7_cond <= VAR_t8_MUX_uxn_opcodes_h_l1809_c2_bab7_cond;
     t8_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue;
     t8_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output := t8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1825_c7_f7c3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output := result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1822_c7_d6d6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_f7c3_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1822_c7_d6d6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output := result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output;

     -- n8_MUX[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1809_c2_bab7_cond <= VAR_n8_MUX_uxn_opcodes_h_l1809_c2_bab7_cond;
     n8_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue;
     n8_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output := n8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_d6d6_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1809_c2_bab7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output := result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1837_l1805_DUPLICATE_6ea5 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1837_l1805_DUPLICATE_6ea5_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_922a(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_bab7_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1837_l1805_DUPLICATE_6ea5_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1837_l1805_DUPLICATE_6ea5_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
