-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 36
entity nip2_0CLK_1a2ef46d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_1a2ef46d;
architecture arch of nip2_0CLK_1a2ef46d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2175_c6_1f5f]
signal BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2175_c2_556d]
signal t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2175_c2_556d]
signal t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2175_c2_556d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2175_c2_556d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2175_c2_556d]
signal result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2175_c2_556d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2175_c2_556d]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2175_c2_556d]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2175_c2_556d]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2175_c2_556d]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2175_c2_556d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2188_c11_c48a]
signal BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2188_c7_0379]
signal t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2188_c7_0379]
signal t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2188_c7_0379]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2188_c7_0379]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2188_c7_0379]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2188_c7_0379]
signal result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2188_c7_0379]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2191_c11_d783]
signal BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2191_c7_7b3c]
signal t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2191_c7_7b3c]
signal t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2191_c7_7b3c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2191_c7_7b3c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2191_c7_7b3c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2191_c7_7b3c]
signal result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2191_c7_7b3c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2193_c30_442b]
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2198_c11_fbad]
signal BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2198_c7_97af]
signal t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2198_c7_97af]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2198_c7_97af]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2198_c7_97af]
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2198_c7_97af]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_return_output : unsigned(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a6df( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_vram_write := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f
BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_left,
BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_right,
BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2175_c2_556d
t16_low_MUX_uxn_opcodes_h_l2175_c2_556d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_cond,
t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue,
t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse,
t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2175_c2_556d
t16_high_MUX_uxn_opcodes_h_l2175_c2_556d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_cond,
t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue,
t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse,
t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_left,
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_right,
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2188_c7_0379
t16_low_MUX_uxn_opcodes_h_l2188_c7_0379 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_cond,
t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue,
t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse,
t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2188_c7_0379
t16_high_MUX_uxn_opcodes_h_l2188_c7_0379 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_cond,
t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue,
t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse,
t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_cond,
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783
BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_left,
BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_right,
BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c
t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond,
t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue,
t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse,
t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c
t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond,
t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue,
t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse,
t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2193_c30_442b
sp_relative_shift_uxn_opcodes_h_l2193_c30_442b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_ins,
sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_x,
sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_y,
sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_left,
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_right,
BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2198_c7_97af
t16_low_MUX_uxn_opcodes_h_l2198_c7_97af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_cond,
t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue,
t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse,
t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_cond,
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output,
 t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
 t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_return_output,
 t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_return_output,
 t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_return_output,
 t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output,
 t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output,
 sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_return_output,
 t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2180_c3_f299 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_9dbb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2189_c3_58cd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2195_c3_37fa : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2200_c3_d876 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2201_c3_a5fe : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2198_c7_97af_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2198_l2188_l2175_DUPLICATE_1faa_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_7145_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2198_l2188_l2191_DUPLICATE_0870_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2191_DUPLICATE_38e4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2206_l2171_DUPLICATE_22a6_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_right := to_unsigned(3, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2201_c3_a5fe := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2201_c3_a5fe;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2180_c3_f299 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2180_c3_f299;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_9dbb := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_9dbb;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2200_c3_d876 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2200_c3_d876;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2195_c3_37fa := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2195_c3_37fa;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2189_c3_58cd := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2189_c3_58cd;
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse := t16_high;
     VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse := t16_low;
     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2175_c2_556d_return_output := result.is_vram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_7145 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_7145_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2198_c11_fbad] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_left;
     BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_return_output := BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2175_c2_556d_return_output := result.is_pc_updated;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2175_c2_556d_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2188_c11_c48a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2193_c30_442b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_ins;
     sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_x;
     sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_return_output := sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2191_c11_d783] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_left;
     BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_return_output := BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2198_c7_97af] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2198_c7_97af_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2198_l2188_l2175_DUPLICATE_1faa LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2198_l2188_l2175_DUPLICATE_1faa_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2191_DUPLICATE_38e4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2191_DUPLICATE_38e4_return_output := result.is_stack_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2175_c2_556d_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2198_l2188_l2191_DUPLICATE_0870 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2198_l2188_l2191_DUPLICATE_0870_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2175_c6_1f5f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2175_c6_1f5f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_c48a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2191_c11_d783_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2198_c11_fbad_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_7145_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2198_l2188_DUPLICATE_7145_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2198_l2188_l2191_DUPLICATE_0870_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2198_l2188_l2191_DUPLICATE_0870_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2198_l2188_l2191_DUPLICATE_0870_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2191_DUPLICATE_38e4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2191_DUPLICATE_38e4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2198_l2188_l2175_DUPLICATE_1faa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2198_l2188_l2175_DUPLICATE_1faa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2198_l2188_l2175_DUPLICATE_1faa_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2175_c2_556d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2175_c2_556d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2175_c2_556d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2175_c2_556d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2198_c7_97af_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_442b_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2198_c7_97af] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_return_output := result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2191_c7_7b3c] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond;
     t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output := t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2191_c7_7b3c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2198_c7_97af] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2198_c7_97af] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2198_c7_97af] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_cond;
     t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_return_output := t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2198_c7_97af] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2198_c7_97af_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2198_c7_97af_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2198_c7_97af_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2198_c7_97af_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2198_c7_97af_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2188_c7_0379] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2191_c7_7b3c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2191_c7_7b3c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2191_c7_7b3c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2188_c7_0379] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_cond;
     t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_return_output := t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2191_c7_7b3c] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond;
     t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output := t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2191_c7_7b3c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2191_c7_7b3c_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2188_c7_0379] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_return_output := result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_cond;
     t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_return_output := t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2188_c7_0379] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2188_c7_0379] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_cond;
     t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_return_output := t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2188_c7_0379] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2188_c7_0379] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2175_c2_556d_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2188_c7_0379_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2175_c2_556d] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_cond;
     t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_return_output := t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_return_output;

     -- Submodule level 5
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2175_c2_556d_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2206_l2171_DUPLICATE_22a6 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2206_l2171_DUPLICATE_22a6_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a6df(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2175_c2_556d_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2206_l2171_DUPLICATE_22a6_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2206_l2171_DUPLICATE_22a6_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
