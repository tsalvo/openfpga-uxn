-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity eor_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor_0CLK_64d180f1;
architecture arch of eor_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1099_c6_22ed]
signal BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1099_c2_7d4f]
signal t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1099_c2_7d4f]
signal n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1099_c2_7d4f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1099_c2_7d4f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1099_c2_7d4f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1099_c2_7d4f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1099_c2_7d4f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1099_c2_7d4f]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1099_c2_7d4f]
signal result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1099_c2_7d4f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1099_c2_7d4f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1112_c11_9e58]
signal BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1112_c7_083a]
signal t8_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1112_c7_083a]
signal n8_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1112_c7_083a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1112_c7_083a]
signal result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1112_c7_083a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1112_c7_083a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1112_c7_083a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1115_c11_7532]
signal BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1115_c7_a0a4]
signal t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1115_c7_a0a4]
signal n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1115_c7_a0a4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1115_c7_a0a4]
signal result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1115_c7_a0a4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1115_c7_a0a4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1115_c7_a0a4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1118_c11_d62e]
signal BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1118_c7_58bc]
signal n8_MUX_uxn_opcodes_h_l1118_c7_58bc_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1118_c7_58bc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1118_c7_58bc]
signal result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1118_c7_58bc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1118_c7_58bc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1118_c7_58bc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1120_c30_f2fd]
signal sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_return_output : signed(3 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1123_c21_edd7]
signal BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_left : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_right : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed
BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_left,
BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_right,
BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output);

-- t8_MUX_uxn_opcodes_h_l1099_c2_7d4f
t8_MUX_uxn_opcodes_h_l1099_c2_7d4f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond,
t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue,
t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse,
t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output);

-- n8_MUX_uxn_opcodes_h_l1099_c2_7d4f
n8_MUX_uxn_opcodes_h_l1099_c2_7d4f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond,
n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue,
n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse,
n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f
result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f
result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f
result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f
result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f
result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f
result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58
BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_left,
BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_right,
BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_return_output);

-- t8_MUX_uxn_opcodes_h_l1112_c7_083a
t8_MUX_uxn_opcodes_h_l1112_c7_083a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1112_c7_083a_cond,
t8_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue,
t8_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse,
t8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output);

-- n8_MUX_uxn_opcodes_h_l1112_c7_083a
n8_MUX_uxn_opcodes_h_l1112_c7_083a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1112_c7_083a_cond,
n8_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue,
n8_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse,
n8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532
BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_left,
BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_right,
BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_return_output);

-- t8_MUX_uxn_opcodes_h_l1115_c7_a0a4
t8_MUX_uxn_opcodes_h_l1115_c7_a0a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond,
t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue,
t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse,
t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output);

-- n8_MUX_uxn_opcodes_h_l1115_c7_a0a4
n8_MUX_uxn_opcodes_h_l1115_c7_a0a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond,
n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue,
n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse,
n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4
result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4
result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4
result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e
BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_left,
BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_right,
BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_return_output);

-- n8_MUX_uxn_opcodes_h_l1118_c7_58bc
n8_MUX_uxn_opcodes_h_l1118_c7_58bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1118_c7_58bc_cond,
n8_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue,
n8_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse,
n8_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc
result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc
result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_cond,
result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc
result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc
result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd
sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_ins,
sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_x,
sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_y,
sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7
BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7 : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_left,
BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_right,
BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output,
 t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
 n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_return_output,
 t8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output,
 n8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_return_output,
 t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output,
 n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_return_output,
 n8_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output,
 sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1104_c3_5bd4 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1109_c3_da4d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1113_c3_a5cd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1118_c7_58bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1122_c3_13e6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_f3c9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_6aae_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_1081_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_1da6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1118_l1115_DUPLICATE_a6ad_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1127_l1095_DUPLICATE_b65c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1122_c3_13e6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1122_c3_13e6;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1109_c3_da4d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1109_c3_da4d;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1113_c3_a5cd := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1113_c3_a5cd;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_right := to_unsigned(2, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_right := to_unsigned(3, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1104_c3_5bd4 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1104_c3_5bd4;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_1da6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_1da6_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1112_c11_9e58] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_left;
     BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_return_output := BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_1081 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_1081_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1099_c6_22ed] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_left;
     BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output := BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output;

     -- BIN_OP_XOR[uxn_opcodes_h_l1123_c21_edd7] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_left;
     BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_return_output := BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1118_l1115_DUPLICATE_a6ad LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1118_l1115_DUPLICATE_a6ad_return_output := result.stack_address_sp_offset;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1099_c2_7d4f_return_output := result.is_ram_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1099_c2_7d4f_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1118_c11_d62e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_f3c9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_f3c9_return_output := result.u8_value;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1099_c2_7d4f_return_output := result.is_pc_updated;

     -- sp_relative_shift[uxn_opcodes_h_l1120_c30_f2fd] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_ins;
     sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_x;
     sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_return_output := sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1099_c2_7d4f_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1115_c11_7532] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_left;
     BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_return_output := BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_6aae LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_6aae_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_22ed_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1112_c7_083a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1112_c7_083a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9e58_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_7532_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1118_c7_58bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_d62e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_edd7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_1081_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_1081_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_1081_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_6aae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_6aae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_6aae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_1da6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_1da6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_1da6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1118_l1115_DUPLICATE_a6ad_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1118_l1115_DUPLICATE_a6ad_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_f3c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_f3c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_f3c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_f3c9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1099_c2_7d4f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1099_c2_7d4f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1099_c2_7d4f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1099_c2_7d4f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_f2fd_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1118_c7_58bc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output := result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1118_c7_58bc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1118_c7_58bc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output;

     -- t8_MUX[uxn_opcodes_h_l1115_c7_a0a4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond <= VAR_t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond;
     t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue;
     t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output := t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1118_c7_58bc] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1118_c7_58bc_cond <= VAR_n8_MUX_uxn_opcodes_h_l1118_c7_58bc_cond;
     n8_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue;
     n8_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output := n8_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1118_c7_58bc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1118_c7_58bc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_58bc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;
     -- t8_MUX[uxn_opcodes_h_l1112_c7_083a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1112_c7_083a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1112_c7_083a_cond;
     t8_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue;
     t8_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output := t8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1115_c7_a0a4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1115_c7_a0a4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1115_c7_a0a4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1115_c7_a0a4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1115_c7_a0a4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond <= VAR_n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond;
     n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue;
     n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output := n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1115_c7_a0a4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_a0a4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;
     -- t8_MUX[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond;
     t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue;
     t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output := t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output;

     -- n8_MUX[uxn_opcodes_h_l1112_c7_083a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1112_c7_083a_cond <= VAR_n8_MUX_uxn_opcodes_h_l1112_c7_083a_cond;
     n8_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue;
     n8_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output := n8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1112_c7_083a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1112_c7_083a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1112_c7_083a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1112_c7_083a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1112_c7_083a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_083a_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output;

     -- n8_MUX[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond;
     n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue;
     n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output := n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1099_c2_7d4f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1127_l1095_DUPLICATE_b65c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1127_l1095_DUPLICATE_b65c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_7d4f_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1127_l1095_DUPLICATE_b65c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1127_l1095_DUPLICATE_b65c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
