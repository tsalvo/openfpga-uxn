-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 55
entity lit_0CLK_3220bbf1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lit_0CLK_3220bbf1;
architecture arch of lit_0CLK_3220bbf1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l206_c6_2572]
signal BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l206_c1_485a]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l206_c2_b3f4]
signal tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l206_c2_b3f4]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l206_c2_b3f4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : signed(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l206_c2_b3f4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(0 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l206_c2_b3f4]
signal result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l206_c2_b3f4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l206_c2_b3f4]
signal result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(7 downto 0);

-- result_is_ram_read_MUX[uxn_opcodes_h_l206_c2_b3f4]
signal result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l206_c2_b3f4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l206_c2_b3f4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l206_c2_b3f4]
signal result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l207_c3_f36b[uxn_opcodes_h_l207_c3_f36b]
signal printf_uxn_opcodes_h_l207_c3_f36b_uxn_opcodes_h_l207_c3_f36b_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l212_c11_635d]
signal BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l212_c7_ad27]
signal tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l212_c7_ad27]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l212_c7_ad27]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(0 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l212_c7_ad27]
signal result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l212_c7_ad27]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l212_c7_ad27]
signal result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(7 downto 0);

-- result_is_ram_read_MUX[uxn_opcodes_h_l212_c7_ad27]
signal result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l212_c7_ad27]
signal result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l212_c7_ad27]
signal result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l212_c7_ad27]
signal result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l217_c11_aef5]
signal BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l217_c7_eb25]
signal tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l217_c7_eb25]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(0 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l217_c7_eb25]
signal result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l217_c7_eb25]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l217_c7_eb25]
signal result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(7 downto 0);

-- result_is_ram_read_MUX[uxn_opcodes_h_l217_c7_eb25]
signal result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l217_c7_eb25]
signal result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l217_c7_eb25]
signal result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l217_c7_eb25]
signal result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l220_c11_f704]
signal BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l220_c7_41af]
signal tmp8_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l220_c7_41af]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l220_c7_41af]
signal result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l220_c7_41af]
signal result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(0 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l220_c7_41af]
signal result_pc_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l220_c7_41af]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l220_c7_41af]
signal result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(7 downto 0);

-- result_is_ram_read_MUX[uxn_opcodes_h_l220_c7_41af]
signal result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l224_c15_6df5]
signal BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l226_c11_0a4f]
signal BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l226_c7_646d]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l226_c7_646d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l226_c7_646d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l226_c7_646d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l226_c7_646d]
signal result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l232_c11_96ac]
signal BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l232_c7_fc04]
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l232_c7_fc04]
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_170c( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : signed;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.sp_relative_shift := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.pc := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.stack_value := ref_toks_6;
      base.is_ram_read := ref_toks_7;
      base.is_stack_write := ref_toks_8;
      base.is_opc_done := ref_toks_9;
      base.ram_addr := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572
BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_left,
BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_right,
BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_return_output);

-- tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4
tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_cond,
tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue,
tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse,
tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4
result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4
result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4
result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output);

-- result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4
result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_cond,
result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue,
result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse,
result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4
result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_cond,
result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output);

-- result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4
result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_cond,
result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue,
result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse,
result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4
result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4
result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4
result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_cond,
result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output);

-- printf_uxn_opcodes_h_l207_c3_f36b_uxn_opcodes_h_l207_c3_f36b
printf_uxn_opcodes_h_l207_c3_f36b_uxn_opcodes_h_l207_c3_f36b : entity work.printf_uxn_opcodes_h_l207_c3_f36b_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l207_c3_f36b_uxn_opcodes_h_l207_c3_f36b_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d
BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_left,
BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_right,
BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output);

-- tmp8_MUX_uxn_opcodes_h_l212_c7_ad27
tmp8_MUX_uxn_opcodes_h_l212_c7_ad27 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_cond,
tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue,
tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse,
tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27
result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27
result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_return_output);

-- result_pc_MUX_uxn_opcodes_h_l212_c7_ad27
result_pc_MUX_uxn_opcodes_h_l212_c7_ad27 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_cond,
result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue,
result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse,
result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27
result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_cond,
result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_return_output);

-- result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27
result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_cond,
result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue,
result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse,
result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27
result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27
result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27
result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_cond,
result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5
BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_left,
BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_right,
BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output);

-- tmp8_MUX_uxn_opcodes_h_l217_c7_eb25
tmp8_MUX_uxn_opcodes_h_l217_c7_eb25 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_cond,
tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue,
tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse,
tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_return_output);

-- result_pc_MUX_uxn_opcodes_h_l217_c7_eb25
result_pc_MUX_uxn_opcodes_h_l217_c7_eb25 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_cond,
result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue,
result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse,
result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25
result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_cond,
result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_return_output);

-- result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25
result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_cond,
result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue,
result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse,
result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25
result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25
result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25
result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_cond,
result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704
BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_left,
BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_right,
BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output);

-- tmp8_MUX_uxn_opcodes_h_l220_c7_41af
tmp8_MUX_uxn_opcodes_h_l220_c7_41af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l220_c7_41af_cond,
tmp8_MUX_uxn_opcodes_h_l220_c7_41af_iftrue,
tmp8_MUX_uxn_opcodes_h_l220_c7_41af_iffalse,
tmp8_MUX_uxn_opcodes_h_l220_c7_41af_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af
result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af
result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af
result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_return_output);

-- result_pc_MUX_uxn_opcodes_h_l220_c7_41af
result_pc_MUX_uxn_opcodes_h_l220_c7_41af : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l220_c7_41af_cond,
result_pc_MUX_uxn_opcodes_h_l220_c7_41af_iftrue,
result_pc_MUX_uxn_opcodes_h_l220_c7_41af_iffalse,
result_pc_MUX_uxn_opcodes_h_l220_c7_41af_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af
result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_cond,
result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_return_output);

-- result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af
result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_cond,
result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_iftrue,
result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_iffalse,
result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5
BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5 : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_left,
BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_right,
BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f
BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_left,
BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_right,
BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d
result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_cond,
result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac
BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_left,
BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_right,
BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_return_output,
 tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
 result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
 result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output,
 tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_return_output,
 result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_return_output,
 result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output,
 tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_return_output,
 result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_return_output,
 result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output,
 tmp8_MUX_uxn_opcodes_h_l220_c7_41af_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_return_output,
 result_pc_MUX_uxn_opcodes_h_l220_c7_41af_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_return_output,
 result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_iffalse : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l209_c3_8cfe : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l206_c2_b3f4_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l207_c3_f36b_uxn_opcodes_h_l207_c3_f36b_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l212_c7_ad27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_uxn_opcodes_h_l224_c3_4e21 : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l229_c3_48aa : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l206_l212_l226_l217_DUPLICATE_f392_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l206_l220_l212_l217_DUPLICATE_da95_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_c20e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_6741_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_read_d41d_uxn_opcodes_h_l206_l220_l217_DUPLICATE_0654_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l217_l212_l206_l232_DUPLICATE_2f2c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l206_l217_DUPLICATE_3419_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l217_l212_l232_l226_DUPLICATE_7729_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_170c_uxn_opcodes_h_l237_l201_DUPLICATE_6fba_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_right := to_unsigned(3, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l209_c3_8cfe := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l209_c3_8cfe;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l229_c3_48aa := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l229_c3_48aa;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_right := to_unsigned(0, 1);
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_iffalse := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_left := VAR_pc;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue := VAR_pc;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_left := VAR_phase;
     VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_41af_iftrue := VAR_previous_ram_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_41af_iffalse := tmp8;
     -- BIN_OP_PLUS[uxn_opcodes_h_l224_c15_6df5] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_left;
     BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_return_output := BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l232_c11_96ac] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_left;
     BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_return_output := BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_read_d41d_uxn_opcodes_h_l206_l220_l217_DUPLICATE_0654 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_read_d41d_uxn_opcodes_h_l206_l220_l217_DUPLICATE_0654_return_output := result.is_ram_read;

     -- result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d[uxn_opcodes_h_l212_c7_ad27] LATENCY=0
     VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l212_c7_ad27_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_c20e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_c20e_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l220_c11_f704] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_left;
     BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output := BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l206_l220_l212_l217_DUPLICATE_da95 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l206_l220_l212_l217_DUPLICATE_da95_return_output := result.pc;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l217_l212_l232_l226_DUPLICATE_7729 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l217_l212_l232_l226_DUPLICATE_7729_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l206_l212_l226_l217_DUPLICATE_f392 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l206_l212_l226_l217_DUPLICATE_f392_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l226_c11_0a4f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_left;
     BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_return_output := BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l217_l212_l206_l232_DUPLICATE_2f2c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l217_l212_l206_l232_DUPLICATE_2f2c_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l206_c6_2572] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_left;
     BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output := BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_6741 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_6741_return_output := result.stack_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l217_c11_aef5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_left;
     BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output := BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l206_l217_DUPLICATE_3419 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l206_l217_DUPLICATE_3419_return_output := result.ram_addr;

     -- BIN_OP_EQ[uxn_opcodes_h_l212_c11_635d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_left;
     BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output := BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l206_c2_b3f4] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l206_c2_b3f4_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_2572_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_635d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_aef5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_41af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_41af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_f704_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_0a4f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_96ac_return_output;
     VAR_result_pc_uxn_opcodes_h_l224_c3_4e21 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_6df5_return_output, 16);
     VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l206_l220_l212_l217_DUPLICATE_da95_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l206_l220_l212_l217_DUPLICATE_da95_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l206_l220_l212_l217_DUPLICATE_da95_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_41af_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l206_l220_l212_l217_DUPLICATE_da95_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l206_l217_DUPLICATE_3419_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l206_l217_DUPLICATE_3419_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l217_l212_l232_l226_DUPLICATE_7729_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l217_l212_l232_l226_DUPLICATE_7729_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l217_l212_l232_l226_DUPLICATE_7729_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l217_l212_l232_l226_DUPLICATE_7729_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l217_l212_l232_l226_DUPLICATE_7729_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l206_l212_l226_l217_DUPLICATE_f392_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l206_l212_l226_l217_DUPLICATE_f392_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l206_l212_l226_l217_DUPLICATE_f392_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l206_l212_l226_l217_DUPLICATE_f392_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_read_d41d_uxn_opcodes_h_l206_l220_l217_DUPLICATE_0654_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_read_d41d_uxn_opcodes_h_l206_l220_l217_DUPLICATE_0654_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_read_d41d_uxn_opcodes_h_l206_l220_l217_DUPLICATE_0654_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l217_l212_l206_l232_DUPLICATE_2f2c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l217_l212_l206_l232_DUPLICATE_2f2c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l217_l212_l206_l232_DUPLICATE_2f2c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l217_l212_l206_l232_DUPLICATE_2f2c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l217_l212_l206_l232_DUPLICATE_2f2c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_c20e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_c20e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_c20e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_c20e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_c20e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_6741_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_6741_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_6741_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_6741_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l217_l212_l206_l226_DUPLICATE_6741_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse := VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l212_c7_ad27_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l206_c2_b3f4_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_41af_iftrue := VAR_result_pc_uxn_opcodes_h_l224_c3_4e21;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l212_c7_ad27] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l220_c7_41af] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l220_c7_41af_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_41af_cond;
     tmp8_MUX_uxn_opcodes_h_l220_c7_41af_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_41af_iftrue;
     tmp8_MUX_uxn_opcodes_h_l220_c7_41af_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_41af_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_41af_return_output := tmp8_MUX_uxn_opcodes_h_l220_c7_41af_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l217_c7_eb25] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_return_output := result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l232_c7_fc04] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l226_c7_646d] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_cond;
     result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_return_output := result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l232_c7_fc04] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l220_c7_41af] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l220_c7_41af_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_41af_cond;
     result_pc_MUX_uxn_opcodes_h_l220_c7_41af_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_41af_iftrue;
     result_pc_MUX_uxn_opcodes_h_l220_c7_41af_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_41af_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_41af_return_output := result_pc_MUX_uxn_opcodes_h_l220_c7_41af_return_output;

     -- result_is_ram_read_MUX[uxn_opcodes_h_l220_c7_41af] LATENCY=0
     -- Inputs
     result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_cond <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_cond;
     result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_iftrue <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_iftrue;
     result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_iffalse <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_iffalse;
     -- Outputs
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_return_output := result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l226_c7_646d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l226_c7_646d] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l206_c1_485a] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l206_c2_b3f4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l207_c3_f36b_uxn_opcodes_h_l207_c3_f36b_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_485a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fc04_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_646d_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse := VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_41af_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fc04_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_41af_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse := VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_646d_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_646d_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_41af_return_output;
     -- result_pc_MUX[uxn_opcodes_h_l217_c7_eb25] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_cond;
     result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue;
     result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_return_output := result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l212_c7_ad27] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_return_output := result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l220_c7_41af] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l220_c7_41af] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_cond;
     result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_return_output := result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l220_c7_41af] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l226_c7_646d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_return_output;

     -- result_is_ram_read_MUX[uxn_opcodes_h_l217_c7_eb25] LATENCY=0
     -- Inputs
     result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_cond <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_cond;
     result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue;
     result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse;
     -- Outputs
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_return_output := result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;

     -- printf_uxn_opcodes_h_l207_c3_f36b[uxn_opcodes_h_l207_c3_f36b] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l207_c3_f36b_uxn_opcodes_h_l207_c3_f36b_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l207_c3_f36b_uxn_opcodes_h_l207_c3_f36b_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_opc_done_MUX[uxn_opcodes_h_l226_c7_646d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l206_c2_b3f4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l217_c7_eb25] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_cond;
     tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue;
     tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_return_output := tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_646d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_41af_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse := VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_646d_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse := VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_41af_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_41af_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l220_c7_41af] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l212_c7_ad27] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_cond;
     tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue;
     tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_return_output := tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l206_c2_b3f4] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output := result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l220_c7_41af] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_return_output;

     -- result_is_ram_read_MUX[uxn_opcodes_h_l212_c7_ad27] LATENCY=0
     -- Inputs
     result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_cond <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_cond;
     result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue;
     result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse;
     -- Outputs
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_return_output := result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l217_c7_eb25] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_cond;
     result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_return_output := result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l217_c7_eb25] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l217_c7_eb25] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l212_c7_ad27] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_cond;
     result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue;
     result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_return_output := result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_41af_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse := VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_41af_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;
     -- result_is_ram_read_MUX[uxn_opcodes_h_l206_c2_b3f4] LATENCY=0
     -- Inputs
     result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_cond <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_cond;
     result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue;
     result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse;
     -- Outputs
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output := result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l212_c7_ad27] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l212_c7_ad27] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l206_c2_b3f4] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_cond;
     result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue;
     result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output := result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l212_c7_ad27] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_cond;
     result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_return_output := result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l217_c7_eb25] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l217_c7_eb25] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l206_c2_b3f4] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_cond;
     tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue;
     tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output := tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_eb25_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l206_c2_b3f4] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l212_c7_ad27] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l206_c2_b3f4] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_cond;
     result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output := result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l212_c7_ad27] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l206_c2_b3f4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_ad27_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l206_c2_b3f4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l206_c2_b3f4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_170c_uxn_opcodes_h_l237_l201_DUPLICATE_6fba LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_170c_uxn_opcodes_h_l237_l201_DUPLICATE_6fba_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_170c(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
     VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output,
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_b3f4_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_170c_uxn_opcodes_h_l237_l201_DUPLICATE_6fba_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_170c_uxn_opcodes_h_l237_l201_DUPLICATE_6fba_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
