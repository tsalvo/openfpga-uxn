-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sth2_0CLK_55b6500a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth2_0CLK_55b6500a;
architecture arch of sth2_0CLK_55b6500a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2419_c6_d33c]
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2419_c2_abfe]
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2419_c2_abfe]
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2419_c2_abfe]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2419_c2_abfe]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2419_c2_abfe]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2419_c2_abfe]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2419_c2_abfe]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2419_c2_abfe]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2419_c2_abfe]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2419_c2_abfe]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2419_c2_abfe]
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2432_c11_7698]
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2432_c7_4768]
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2432_c7_4768]
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2432_c7_4768]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2432_c7_4768]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2432_c7_4768]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2432_c7_4768]
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2432_c7_4768]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2432_c7_4768]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2435_c11_f633]
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2435_c7_84cf]
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2435_c7_84cf]
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2435_c7_84cf]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2435_c7_84cf]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2435_c7_84cf]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2435_c7_84cf]
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2435_c7_84cf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2435_c7_84cf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2437_c30_2a5d]
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2439_c11_2eaa]
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2439_c7_b4e7]
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2439_c7_b4e7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2439_c7_b4e7]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2439_c7_b4e7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2439_c7_b4e7]
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2439_c7_b4e7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2439_c7_b4e7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2447_c11_c2bc]
signal BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2447_c7_0b62]
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2447_c7_0b62]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2447_c7_0b62]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2447_c7_0b62]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8b52( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_left,
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_right,
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe
t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_cond,
t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue,
t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse,
t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe
t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_cond,
t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue,
t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse,
t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_cond,
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_left,
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_right,
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2432_c7_4768
t16_low_MUX_uxn_opcodes_h_l2432_c7_4768 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_cond,
t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue,
t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse,
t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2432_c7_4768
t16_high_MUX_uxn_opcodes_h_l2432_c7_4768 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_cond,
t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue,
t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse,
t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_cond,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_left,
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_right,
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf
t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_cond,
t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue,
t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse,
t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf
t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_cond,
t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue,
t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse,
t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_cond,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d
sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_ins,
sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_x,
sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_y,
sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_left,
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_right,
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7
t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond,
t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue,
t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse,
t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond,
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_left,
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_right,
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_cond,
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output,
 t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
 t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output,
 t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_return_output,
 t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output,
 t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output,
 t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output,
 sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_return_output,
 t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2424_c3_5330 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_c7d7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_9d06 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2442_c3_fbab : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2444_c3_8d68 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2448_c3_ab50 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2449_c3_a70b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_342d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_a293_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_886b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_e5ed_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_300a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_968d_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2454_l2415_DUPLICATE_f2dc_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_y := resize(to_signed(-2, 3), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_c7d7 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_c7d7;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2424_c3_5330 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2424_c3_5330;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_9d06 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_9d06;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2442_c3_fbab := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2442_c3_fbab;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2449_c3_a70b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2449_c3_a70b;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2444_c3_8d68 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2444_c3_8d68;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2448_c3_ab50 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2448_c3_ab50;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_left := VAR_phase;
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse := t16_high;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse := t16_low;
     -- BIN_OP_EQ[uxn_opcodes_h_l2447_c11_c2bc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_left;
     BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_return_output := BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2419_c2_abfe_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_968d LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_968d_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l2437_c30_2a5d] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_ins;
     sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_x;
     sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_return_output := sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2419_c2_abfe_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2432_c11_7698] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_left;
     BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output := BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_886b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_886b_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2419_c6_d33c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2419_c2_abfe_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2435_c11_f633] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_left;
     BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output := BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2439_c11_2eaa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_left;
     BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_return_output := BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_a293 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_a293_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_300a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_300a_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_342d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_342d_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_e5ed LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_e5ed_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_d33c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_7698_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_f633_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2eaa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_c2bc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_a293_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_a293_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_300a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_300a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_300a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_300a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_886b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_886b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_886b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_e5ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_e5ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_e5ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_968d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_968d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_342d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_342d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_342d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_342d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2419_c2_abfe_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2419_c2_abfe_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2419_c2_abfe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_2a5d_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2447_c7_0b62] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2447_c7_0b62] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2435_c7_84cf] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_cond;
     t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output := t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2447_c7_0b62] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output := result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2439_c7_b4e7] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2439_c7_b4e7] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond;
     t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output := t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2447_c7_0b62] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2439_c7_b4e7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_0b62_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2439_c7_b4e7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2439_c7_b4e7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2435_c7_84cf] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2439_c7_b4e7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2435_c7_84cf] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_cond;
     t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output := t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2439_c7_b4e7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output := result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2432_c7_4768] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_cond;
     t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_return_output := t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2435_c7_84cf] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_b4e7_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2432_c7_4768] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2432_c7_4768] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_cond;
     t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_return_output := t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2432_c7_4768] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2435_c7_84cf] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output := result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2435_c7_84cf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2435_c7_84cf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2435_c7_84cf] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_cond;
     t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output := t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_84cf_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2432_c7_4768] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_return_output := result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_cond;
     t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output := t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2432_c7_4768] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2432_c7_4768] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2432_c7_4768] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_4768_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2419_c2_abfe] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output := result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2454_l2415_DUPLICATE_f2dc LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2454_l2415_DUPLICATE_f2dc_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8b52(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_abfe_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2454_l2415_DUPLICATE_f2dc_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2454_l2415_DUPLICATE_f2dc_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
