-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity gth_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end gth_0CLK_226c8821;
architecture arch of gth_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1827_c6_3a6d]
signal BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1827_c2_b60e]
signal t8_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1827_c2_b60e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1827_c2_b60e]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1827_c2_b60e]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1827_c2_b60e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1827_c2_b60e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1827_c2_b60e]
signal result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1827_c2_b60e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1827_c2_b60e]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1827_c2_b60e]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1827_c2_b60e]
signal n8_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1840_c11_8f1b]
signal BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1840_c7_06b6]
signal t8_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1840_c7_06b6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1840_c7_06b6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1840_c7_06b6]
signal result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1840_c7_06b6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1840_c7_06b6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1840_c7_06b6]
signal n8_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1843_c11_b96a]
signal BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1843_c7_8b00]
signal t8_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1843_c7_8b00]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1843_c7_8b00]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1843_c7_8b00]
signal result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1843_c7_8b00]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1843_c7_8b00]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1843_c7_8b00]
signal n8_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1846_c11_8821]
signal BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1846_c7_3d98]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1846_c7_3d98]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1846_c7_3d98]
signal result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1846_c7_3d98]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1846_c7_3d98]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1846_c7_3d98]
signal n8_MUX_uxn_opcodes_h_l1846_c7_3d98_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1848_c30_ec79]
signal sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_return_output : signed(3 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1851_c21_d0fb]
signal BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_right : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1851_c21_7c0a]
signal MUX_uxn_opcodes_h_l1851_c21_7c0a_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1851_c21_7c0a_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1851_c21_7c0a_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1851_c21_7c0a_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c580( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.u8_value := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d
BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_left,
BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_right,
BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output);

-- t8_MUX_uxn_opcodes_h_l1827_c2_b60e
t8_MUX_uxn_opcodes_h_l1827_c2_b60e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1827_c2_b60e_cond,
t8_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue,
t8_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse,
t8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e
result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e
result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e
result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e
result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e
result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e
result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output);

-- n8_MUX_uxn_opcodes_h_l1827_c2_b60e
n8_MUX_uxn_opcodes_h_l1827_c2_b60e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1827_c2_b60e_cond,
n8_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue,
n8_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse,
n8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b
BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_left,
BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_right,
BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_return_output);

-- t8_MUX_uxn_opcodes_h_l1840_c7_06b6
t8_MUX_uxn_opcodes_h_l1840_c7_06b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1840_c7_06b6_cond,
t8_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue,
t8_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse,
t8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6
result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6
result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_cond,
result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6
result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6
result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output);

-- n8_MUX_uxn_opcodes_h_l1840_c7_06b6
n8_MUX_uxn_opcodes_h_l1840_c7_06b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1840_c7_06b6_cond,
n8_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue,
n8_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse,
n8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a
BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_left,
BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_right,
BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_return_output);

-- t8_MUX_uxn_opcodes_h_l1843_c7_8b00
t8_MUX_uxn_opcodes_h_l1843_c7_8b00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1843_c7_8b00_cond,
t8_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue,
t8_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse,
t8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00
result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00
result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_cond,
result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00
result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00
result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output);

-- n8_MUX_uxn_opcodes_h_l1843_c7_8b00
n8_MUX_uxn_opcodes_h_l1843_c7_8b00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1843_c7_8b00_cond,
n8_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue,
n8_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse,
n8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821
BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_left,
BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_right,
BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98
result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98
result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_cond,
result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98
result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98
result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output);

-- n8_MUX_uxn_opcodes_h_l1846_c7_3d98
n8_MUX_uxn_opcodes_h_l1846_c7_3d98 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1846_c7_3d98_cond,
n8_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue,
n8_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse,
n8_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79
sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_ins,
sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_x,
sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_y,
sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb
BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb : entity work.BIN_OP_GT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_left,
BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_right,
BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_return_output);

-- MUX_uxn_opcodes_h_l1851_c21_7c0a
MUX_uxn_opcodes_h_l1851_c21_7c0a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1851_c21_7c0a_cond,
MUX_uxn_opcodes_h_l1851_c21_7c0a_iftrue,
MUX_uxn_opcodes_h_l1851_c21_7c0a_iffalse,
MUX_uxn_opcodes_h_l1851_c21_7c0a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output,
 t8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
 n8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_return_output,
 t8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output,
 n8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_return_output,
 t8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output,
 n8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output,
 n8_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output,
 sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_return_output,
 MUX_uxn_opcodes_h_l1851_c21_7c0a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1837_c3_b003 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1832_c3_1a76 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1827_c2_b60e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1841_c3_5c6f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1840_c7_06b6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1843_c7_8b00_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1850_c3_3143 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1846_c7_3d98_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1851_c21_7c0a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1851_c21_7c0a_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1851_c21_7c0a_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1851_c21_7c0a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1840_l1843_l1827_l1846_DUPLICATE_d62d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_f778_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_f21f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_16d9_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1843_l1846_DUPLICATE_adfa_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l1823_l1855_DUPLICATE_a0d0_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1832_c3_1a76 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1832_c3_1a76;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1850_c3_3143 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1850_c3_3143;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1837_c3_b003 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1837_c3_b003;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_right := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1851_c21_7c0a_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1851_c21_7c0a_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1841_c3_5c6f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1841_c3_5c6f;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_f21f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_f21f_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1846_c11_8821] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_left;
     BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_return_output := BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_16d9 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_16d9_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1843_l1846_DUPLICATE_adfa LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1843_l1846_DUPLICATE_adfa_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1840_l1843_l1827_l1846_DUPLICATE_d62d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1840_l1843_l1827_l1846_DUPLICATE_d62d_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_f778 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_f778_return_output := result.is_opc_done;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1827_c2_b60e_return_output := result.is_vram_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1827_c2_b60e_return_output := result.is_ram_write;

     -- sp_relative_shift[uxn_opcodes_h_l1848_c30_ec79] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_ins;
     sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_x;
     sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_return_output := sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1851_c21_d0fb] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_left;
     BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_return_output := BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1827_c6_3a6d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1827_c2_b60e_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1840_c11_8f1b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1843_c11_b96a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1827_c2_b60e_return_output := result.is_stack_index_flipped;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1827_c2_b60e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1827_c2_b60e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1827_c6_3a6d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1840_c7_06b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1840_c7_06b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1840_c11_8f1b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1843_c7_8b00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1843_c7_8b00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1843_c11_b96a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1846_c7_3d98_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1846_c11_8821_return_output;
     VAR_MUX_uxn_opcodes_h_l1851_c21_7c0a_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1851_c21_d0fb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_16d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_16d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_16d9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_f778_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_f778_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_f778_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_f21f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_f21f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1840_l1843_l1846_DUPLICATE_f21f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1843_l1846_DUPLICATE_adfa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1843_l1846_DUPLICATE_adfa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1840_l1843_l1827_l1846_DUPLICATE_d62d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1840_l1843_l1827_l1846_DUPLICATE_d62d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1840_l1843_l1827_l1846_DUPLICATE_d62d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1840_l1843_l1827_l1846_DUPLICATE_d62d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1827_c2_b60e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1827_c2_b60e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1827_c2_b60e_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1827_c2_b60e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1848_c30_ec79_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1846_c7_3d98] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1846_c7_3d98] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1846_c7_3d98] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1846_c7_3d98] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output;

     -- t8_MUX[uxn_opcodes_h_l1843_c7_8b00] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1843_c7_8b00_cond <= VAR_t8_MUX_uxn_opcodes_h_l1843_c7_8b00_cond;
     t8_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue;
     t8_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output := t8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;

     -- MUX[uxn_opcodes_h_l1851_c21_7c0a] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1851_c21_7c0a_cond <= VAR_MUX_uxn_opcodes_h_l1851_c21_7c0a_cond;
     MUX_uxn_opcodes_h_l1851_c21_7c0a_iftrue <= VAR_MUX_uxn_opcodes_h_l1851_c21_7c0a_iftrue;
     MUX_uxn_opcodes_h_l1851_c21_7c0a_iffalse <= VAR_MUX_uxn_opcodes_h_l1851_c21_7c0a_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1851_c21_7c0a_return_output := MUX_uxn_opcodes_h_l1851_c21_7c0a_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output;

     -- n8_MUX[uxn_opcodes_h_l1846_c7_3d98] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1846_c7_3d98_cond <= VAR_n8_MUX_uxn_opcodes_h_l1846_c7_3d98_cond;
     n8_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue;
     n8_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output := n8_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue := VAR_MUX_uxn_opcodes_h_l1851_c21_7c0a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;
     -- t8_MUX[uxn_opcodes_h_l1840_c7_06b6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1840_c7_06b6_cond <= VAR_t8_MUX_uxn_opcodes_h_l1840_c7_06b6_cond;
     t8_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue;
     t8_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output := t8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1843_c7_8b00] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1843_c7_8b00] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1846_c7_3d98] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output := result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1843_c7_8b00] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1843_c7_8b00] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;

     -- n8_MUX[uxn_opcodes_h_l1843_c7_8b00] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1843_c7_8b00_cond <= VAR_n8_MUX_uxn_opcodes_h_l1843_c7_8b00_cond;
     n8_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue;
     n8_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output := n8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1846_c7_3d98_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1840_c7_06b6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;

     -- t8_MUX[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1827_c2_b60e_cond <= VAR_t8_MUX_uxn_opcodes_h_l1827_c2_b60e_cond;
     t8_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue;
     t8_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output := t8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1843_c7_8b00] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output := result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1840_c7_06b6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;

     -- n8_MUX[uxn_opcodes_h_l1840_c7_06b6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1840_c7_06b6_cond <= VAR_n8_MUX_uxn_opcodes_h_l1840_c7_06b6_cond;
     n8_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue;
     n8_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output := n8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1840_c7_06b6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1840_c7_06b6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1843_c7_8b00_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output;

     -- n8_MUX[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1827_c2_b60e_cond <= VAR_n8_MUX_uxn_opcodes_h_l1827_c2_b60e_cond;
     n8_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue;
     n8_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output := n8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1840_c7_06b6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output := result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1840_c7_06b6_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1827_c2_b60e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l1823_l1855_DUPLICATE_a0d0 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l1823_l1855_DUPLICATE_a0d0_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c580(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1827_c2_b60e_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l1823_l1855_DUPLICATE_a0d0_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l1823_l1855_DUPLICATE_a0d0_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
