-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity lth_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lth_0CLK_226c8821;
architecture arch of lth_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1889_c6_4c66]
signal BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1889_c2_95d8]
signal result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1889_c2_95d8]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1889_c2_95d8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1889_c2_95d8]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1889_c2_95d8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1889_c2_95d8]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1889_c2_95d8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1889_c2_95d8]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1889_c2_95d8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1889_c2_95d8]
signal n8_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1889_c2_95d8]
signal t8_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1902_c11_530b]
signal BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1902_c7_a13f]
signal result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1902_c7_a13f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1902_c7_a13f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1902_c7_a13f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1902_c7_a13f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1902_c7_a13f]
signal n8_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1902_c7_a13f]
signal t8_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1905_c11_35e5]
signal BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1905_c7_0626]
signal result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1905_c7_0626]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1905_c7_0626]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1905_c7_0626]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1905_c7_0626]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1905_c7_0626]
signal n8_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1905_c7_0626]
signal t8_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1908_c11_89ec]
signal BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1908_c7_c6b1]
signal result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1908_c7_c6b1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1908_c7_c6b1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1908_c7_c6b1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1908_c7_c6b1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1908_c7_c6b1]
signal n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1910_c30_d54b]
signal sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_return_output : signed(3 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l1913_c21_9973]
signal BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1913_c21_8968]
signal MUX_uxn_opcodes_h_l1913_c21_8968_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1913_c21_8968_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1913_c21_8968_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1913_c21_8968_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_922a( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_pc_updated := ref_toks_6;
      base.is_opc_done := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66
BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_left,
BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_right,
BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8
result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_cond,
result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8
result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8
result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8
result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8
result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8
result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8
result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output);

-- n8_MUX_uxn_opcodes_h_l1889_c2_95d8
n8_MUX_uxn_opcodes_h_l1889_c2_95d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1889_c2_95d8_cond,
n8_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue,
n8_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse,
n8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output);

-- t8_MUX_uxn_opcodes_h_l1889_c2_95d8
t8_MUX_uxn_opcodes_h_l1889_c2_95d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1889_c2_95d8_cond,
t8_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue,
t8_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse,
t8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b
BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_left,
BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_right,
BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f
result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f
result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f
result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output);

-- n8_MUX_uxn_opcodes_h_l1902_c7_a13f
n8_MUX_uxn_opcodes_h_l1902_c7_a13f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1902_c7_a13f_cond,
n8_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue,
n8_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse,
n8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output);

-- t8_MUX_uxn_opcodes_h_l1902_c7_a13f
t8_MUX_uxn_opcodes_h_l1902_c7_a13f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1902_c7_a13f_cond,
t8_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue,
t8_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse,
t8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5
BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_left,
BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_right,
BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626
result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_cond,
result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626
result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626
result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626
result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_return_output);

-- n8_MUX_uxn_opcodes_h_l1905_c7_0626
n8_MUX_uxn_opcodes_h_l1905_c7_0626 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1905_c7_0626_cond,
n8_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue,
n8_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse,
n8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output);

-- t8_MUX_uxn_opcodes_h_l1905_c7_0626
t8_MUX_uxn_opcodes_h_l1905_c7_0626 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1905_c7_0626_cond,
t8_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue,
t8_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse,
t8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec
BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_left,
BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_right,
BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1
result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond,
result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1
result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1
result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1
result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output);

-- n8_MUX_uxn_opcodes_h_l1908_c7_c6b1
n8_MUX_uxn_opcodes_h_l1908_c7_c6b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond,
n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue,
n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse,
n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b
sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_ins,
sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_x,
sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_y,
sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973
BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973 : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_left,
BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_right,
BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_return_output);

-- MUX_uxn_opcodes_h_l1913_c21_8968
MUX_uxn_opcodes_h_l1913_c21_8968 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1913_c21_8968_cond,
MUX_uxn_opcodes_h_l1913_c21_8968_iftrue,
MUX_uxn_opcodes_h_l1913_c21_8968_iffalse,
MUX_uxn_opcodes_h_l1913_c21_8968_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
 n8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
 t8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output,
 n8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output,
 t8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_return_output,
 n8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output,
 t8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output,
 n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output,
 sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_return_output,
 BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_return_output,
 MUX_uxn_opcodes_h_l1913_c21_8968_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1899_c3_f51f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1894_c3_26ac : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1889_c2_95d8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1903_c3_3288 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1902_c7_a13f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1905_c7_0626_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1912_c3_a23b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1913_c21_8968_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1913_c21_8968_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1913_c21_8968_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1913_c21_8968_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1889_l1908_l1902_l1905_DUPLICATE_ba14_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_eecc_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_409d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_e3ba_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1908_l1905_DUPLICATE_0eff_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1917_l1885_DUPLICATE_b1f2_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_right := to_unsigned(2, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1912_c3_a23b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1912_c3_a23b;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_right := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1913_c21_8968_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1899_c3_f51f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1899_c3_f51f;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1913_c21_8968_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1903_c3_3288 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1903_c3_3288;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1894_c3_26ac := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1894_c3_26ac;
     VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse := t8;
     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1889_c2_95d8_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1889_l1908_l1902_l1905_DUPLICATE_ba14 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1889_l1908_l1902_l1905_DUPLICATE_ba14_return_output := result.u8_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1889_c2_95d8_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_409d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_409d_return_output := result.is_opc_done;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1889_c2_95d8_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_e3ba LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_e3ba_return_output := result.is_stack_write;

     -- BIN_OP_LT[uxn_opcodes_h_l1913_c21_9973] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_left;
     BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_return_output := BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_eecc LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_eecc_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1902_c11_530b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1908_l1905_DUPLICATE_0eff LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1908_l1905_DUPLICATE_0eff_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1889_c2_95d8_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1905_c11_35e5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1910_c30_d54b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_ins;
     sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_x;
     sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_return_output := sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1889_c6_4c66] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_left;
     BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output := BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1908_c11_89ec] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_left;
     BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_return_output := BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1889_c2_95d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1889_c2_95d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1889_c6_4c66_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1902_c7_a13f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1902_c7_a13f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1902_c11_530b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1905_c7_0626_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1905_c7_0626_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1905_c11_35e5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1908_c11_89ec_return_output;
     VAR_MUX_uxn_opcodes_h_l1913_c21_8968_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l1913_c21_9973_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_eecc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_eecc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_eecc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_409d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_409d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_409d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_e3ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_e3ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1908_l1902_l1905_DUPLICATE_e3ba_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1908_l1905_DUPLICATE_0eff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1908_l1905_DUPLICATE_0eff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1889_l1908_l1902_l1905_DUPLICATE_ba14_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1889_l1908_l1902_l1905_DUPLICATE_ba14_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1889_l1908_l1902_l1905_DUPLICATE_ba14_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1889_l1908_l1902_l1905_DUPLICATE_ba14_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1889_c2_95d8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1889_c2_95d8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1889_c2_95d8_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1889_c2_95d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1910_c30_d54b_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1908_c7_c6b1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1908_c7_c6b1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1908_c7_c6b1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output;

     -- n8_MUX[uxn_opcodes_h_l1908_c7_c6b1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond <= VAR_n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond;
     n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue;
     n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output := n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1908_c7_c6b1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output;

     -- MUX[uxn_opcodes_h_l1913_c21_8968] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1913_c21_8968_cond <= VAR_MUX_uxn_opcodes_h_l1913_c21_8968_cond;
     MUX_uxn_opcodes_h_l1913_c21_8968_iftrue <= VAR_MUX_uxn_opcodes_h_l1913_c21_8968_iftrue;
     MUX_uxn_opcodes_h_l1913_c21_8968_iffalse <= VAR_MUX_uxn_opcodes_h_l1913_c21_8968_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1913_c21_8968_return_output := MUX_uxn_opcodes_h_l1913_c21_8968_return_output;

     -- t8_MUX[uxn_opcodes_h_l1905_c7_0626] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1905_c7_0626_cond <= VAR_t8_MUX_uxn_opcodes_h_l1905_c7_0626_cond;
     t8_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue;
     t8_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output := t8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue := VAR_MUX_uxn_opcodes_h_l1913_c21_8968_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;
     -- n8_MUX[uxn_opcodes_h_l1905_c7_0626] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1905_c7_0626_cond <= VAR_n8_MUX_uxn_opcodes_h_l1905_c7_0626_cond;
     n8_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue;
     n8_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output := n8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1905_c7_0626] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1905_c7_0626] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;

     -- t8_MUX[uxn_opcodes_h_l1902_c7_a13f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1902_c7_a13f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1902_c7_a13f_cond;
     t8_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue;
     t8_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output := t8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1905_c7_0626] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1905_c7_0626] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1908_c7_c6b1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output := result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1908_c7_c6b1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1902_c7_a13f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1902_c7_a13f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;

     -- n8_MUX[uxn_opcodes_h_l1902_c7_a13f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1902_c7_a13f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1902_c7_a13f_cond;
     n8_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue;
     n8_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output := n8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1902_c7_a13f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1905_c7_0626] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_return_output := result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1902_c7_a13f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1889_c2_95d8_cond <= VAR_t8_MUX_uxn_opcodes_h_l1889_c2_95d8_cond;
     t8_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue;
     t8_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output := t8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1905_c7_0626_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output;

     -- n8_MUX[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1889_c2_95d8_cond <= VAR_n8_MUX_uxn_opcodes_h_l1889_c2_95d8_cond;
     n8_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue;
     n8_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output := n8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1902_c7_a13f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1902_c7_a13f_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1889_c2_95d8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output := result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1917_l1885_DUPLICATE_b1f2 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1917_l1885_DUPLICATE_b1f2_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_922a(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1889_c2_95d8_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1917_l1885_DUPLICATE_b1f2_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1917_l1885_DUPLICATE_b1f2_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
